��/  {��m݄i�k�ێ]��;�ly�WJ��S���J��S���J��S���J��S���J��S�����&�������nJ��S����㖿UpK�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-�=O ��-���QE����r�����/U�#�k?�M������P:խrQV*��\u�Q�o�����q�<��g:�Bح%�R��2Dp�ݏ~�e�ph9!�4�hԚԾ3�L�AM�G�̴�t�s|B�VT�́:j���+�C`�AF�^ɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<eɽ�*<eɽ�*<e�MO�~I�����1V�@����A�hX@��ω/M|�6��V�!GA>>�-^wq0�	⏌��n~�U���^xω/M|�6��V�!GA>>�-^wq0�Ks�b� �e�`䷟����{v���ԛ��9.[PL�a�X�:霐��{ѧ���9HO��.�vh�F E�L�a�X�:霐��{ѧ���9H`S��|�h.g�/�B�VT�́e���c�t���̌���}O���Nc�T���֤�T�s�D
��[t���̌���}O���Nc�T��w�~Ġ��`��j���f�I�D�J�y�t�h��3����}X|W?+~I�)�]���y���/\�&:�e=AV��3����}X|W?+~I�)�]��wl�=P'���[�I�sʶ��6L����6�c���Z0B��E�I	��o�A�iz�'kL�9�6���귝���Z0B��E�I	��o�A�iz�'k�At����������͗w�)3���jI~�[���@����9��C�'mC�q�X�<QPmssU�*�%-oԕ.���9f?9��C�'mC�q�X�<Q����V
`����]�� �ϵ%[�+ŉ��(l'�<��|����QU��m�q&��a�]mZ�ȟh����iƅ����QU��m�q&���^���$q^�.�2�MuC�l�gd�ѕ�(_:K��.�u��^5�u�,."�9A�F�m �
�\ү�r��M,J�����^5�u�,."�9A�F�m �
�X<Ҹ(ML��2���A`��Cr�A�hX@�������;�,."�9A�F�m �
�\ү�r�z���A��L��{�V�!GA>>�-^wq0�Ks�b� �e�`䷟����{v����W�8��E� ���n�9:霐��{ѧ���9HO��.�vh�F E� ���n�9:霐��{ѧ���9H`S��|�h.g�/�B�VT�́-D�҉%Hj�����x����}O���Nc�T���֤�T�s�D
��[�����x����}O���Nc�T��w�~Ġ��S�Di���{T�_0�����pK�Z���!p=��:霐��{ѧ���9HO��.���Y�1H�愋d�z�}X|W?+~I�)�]��wl�=P'���[�I�sʶ��6L&ꬶ�R\��b�|�� _�5yoɽ�*<eɽ�*<e,4���?wɽ�*<eɽ�*<eɽ�*<e����F�'��zb���<щ��2]|B�~W���J��.�6�o�&�N�`?=ɽ�*<eɽ�*<e�F�:�J�3%7|P�s�%�6ڭWH����	�;�;����-5�M��δ8?Cv.�6�o�&�c�����y�ճ��}�����;��F�t�e����]!�u�"J�ɽ�*<e�VJUT���j+�Xe)����K���L���n�&�G:fGv�A_��l��h�6���δ8?Cvi�OϿY�M�L>�;>c���8��2]|B�~W���J���:eLE7�O��"ɽ�*<eɽ�*<e��2�i;cti�QU�F}nUD�DDHs��G5vb����(�C�I�B?�\���ֻ'�̩;IJvw;ۙ��zN�����>[��H����G:fGv���^�I�ɽ�*<eɽ�*<e����n��r�;&����i��\;�&�����m=b����(�C�I�B?�\���ֻ'i��\;�&y*����i��H�X�I���J��^��k)ɬ׼W��#T�m�2��&�ɽ�*<e��2�i;cti�QU�F�!0K�U&�w�h��t8� @V��	�4�ڟ���u���RΗCf�|��Д�٪,�j�M��gt&ꬶ�R�� �3Y�S���q|���/���?��!f�� �fɽ�*<eC�I k�b����(�C�I�B?�\���ֻ'i��\;�&��z�IYLy��W���S�$o>5����	�;�;���%e�܉<��q��M�ɽ�*<e���J��i�OϿY��,QP��ɽ�*<eɽ�*<e��2�i;cti�QU�FV�v�Ee��V�Q��HO��]��s���RL��F�t�e�7��r|���>�K�R;�e(<�KB\���ֻ'^{�1u$�+���V��.ɽ�*<eɽ�*<e\�@?<�����;.��LQ{D�뫩��[�����K�P ��謋:1.�ez7�i�OϿY�^|��]`�m`�| �s�ڢ>�������K�P ��謋:��9�E"Mc-0��P��T�+Tn��@�7�*,B��z�b�O)ɠo>f�
Y\�er"�꺯z^#w���W����{^�u�P�+H�"�܃$���Zwax8<���3%7|P��LnzI�k����o=/���>;�#���~�ז�t8� @V��	�4�ڟ��o�e�o��T�����)��n�e�j�k�%:Wɓrw�h,*�0�iaɽ�*<e�t8� @V��	�4�ڟ��ʉd��g��g� ���Mh�]=���o�3%7|P��&ʚ�8��F{N.JN{�R�wh�=^f�E���v�"Gs�}�_�av"�v���;�2]|B�~W�t8� @V��	�4�ڟ��ʉd��g��d��w�,�{�`��|�'B������=��>���-5�M�t8� @V��	�4�ڟ�h��1���d��w�,u�P�+H�"�܃$���Zwax8<���3%7|P��LnzI�k�F{N.J��@��MD��`ܖn��t8� @V��	�4�ڟ�h��1��Xz)�aTQT5p`�2|�	R��-L��[��knm`�| �8�1���E������K�P ��謋:�V�旾s�I�`�q��m�2��&��^s�ģ�����^B%4�@_t��ҫ�0�7ӧ�ye�|�	R��-L,��vf�}m`�| �s�ڢ>�������K�P ��謋:�V�旾s�I�`�q�������C��^s�ģ�����^B%4�@_t��ҫ�0�7�i���!�)�2D�5�O㳢mgV�2�OG}Db���q�c�Zwax8<���3%7|P��LnzI�k�����x���8��$����dFK��"Q���X��ViMc�b����(�C�I�B?�Iή�%`���w$o���i��g�����7f6{�~H�@y�����^B%C=֡���)�ߙmit����
���2sdrv��Å����K�P ��謋::a���S�T̨̻v��8<����Iή�%`���[��knm`�| �s�ڢ>�������K�P ��謋:M�TqSݲSAJ��\�~�T�+Tn�iƅ�!8kw��\O)ɠo>f�
Y\�er"�꺯z^ء�s�m.2>���u�P�+H�"�܃$���Zwax8<���3%7|P��LnzI�k7��ɇ�F�/���>;�#���~�ז�t8� @V��	�4�ڟ��y�?=�#,�ry�k���n�e�j���,d�?�����	��,*�0�ia�2]|B�~W�t8� @V��	�4�ڟ���
�(G�y��5����N�`?=|�'B�����\�Co�a3#L�Í����ޞ��K�����N���(����=�/���?��m`�| ��į�O�x�����K�P ��謋:M�TqSݲ�k�UhU�G���2�@k�^s�ģ�����^B%4�@_t���I�\�m�ʱ��
���25��)ϋ�����3�`\\����E�����#~H�@y�����^B%C=֡��͉�+ v����P�6;7}��m4�OO�2ޑ�/���?���V�Q��HO��]��?P�{T���Jnj���hM'��IN��� ��ɢ���2�t8� @V��	�4�ڟ���
�(G�Ɖ�D��0L�O��"�F�:�J�3%7|P��&ʚ�8�t���̌/���>;�#O�bJŤ<�if2>�����] �, ��q�c�Zwax8<���3%7|P��LnzI�k�ϝO�}���8��$������Z0B��l"~<�m	�ViMc�b����(�C�I�B?���3�����w$o���i��g�����7f6{�~H�@y�����^B%C=֡��́��]-�����
���2sdrv��Å����K�P ��謋:x����@j) ����i�8<������3�����[��knm`�| �s�ڢ>�������K�P ��謋:M�TqSݲu�Xn�۸�T�+Tn�iƅ�!�a%�c!O)ɠo>f�
Y\�er"�꺯z^ء�s�m�X�s�Q^�u�P�+H�"�܃$���Zwax8<���3%7|P��LnzI�k(�2Y�ǫ/���>;�#���~�ז�t8� @V��	�4�ڟ��y�?=�#,����N�B��n�e�j���,d�?��i�W��r,*�0�ia�2]|B�~W�t8� @V��	�4�ڟ���
�(G���R���N�`?=|�'B����5>�a��}�a3#L�Í����ޞ��K�����N���(�H���5�/���?��m`�| ��į�O�x�����K�P ��謋:M�TqSݲ��q�6x����2�@k�^s�ģ�����^B%4�@_t��I�b�H汁�
���25��)ϋ�qId�UB\\����E�����#~H�@y�����^B%C=֡���;	��7�8��P�6;7}��m4ک���0[�/���?���V�Q��HO��]��?P�{T��`���$���hM'��IN��� ��ɢ���2�t8� @V��	�4�ڟ���
�(G�r)1�ڹ��O��"�F�:�J�3%7|P��&ʚ�8��s7�}��/���>;�#O�bJŤ<�*��c�P���] �, ��q�c�Zwax8<���3%7|P��LnzI�kdf!п���8��$������Z0B��~,J� ��ViMc�b����(�C�I�B?��x�#αh��w$o���i��g�����7f6{�~H�@y�����^B%C=֡���@w��������
���2sdrv��Å����K�P ��謋:x����@j)�����c^8<�����x�#αh��[��knm`�| �8�1���E������K�P ��謋:�x�A-����Aau�x��j��^s�ģ�����^B%4�@_t���b4?�n"��[�[]��H�(�Ŕ�=�����jt����q�c�Zwax8<���3%7|P��LnzI�kT��82�9��P�6;7}�i�,�N�}74�/���?���V�Q��HO��]��?P�{T�E)�dC��/���?��m`�| ��į�O�x�����K�P ��謋:�x�A-��/���>;�#���7H��^s�ģ�����^B%4�@_t��׷�����0��n�e�j��w��nR>���[��knm`�| �8�1���E������K�P ��謋:�x�A-���ϯ�㳔J�W������^s�ģ�����^B%4�@_t��AC�c�Z�hh�J�.�~-� �����*��I���q�c�Zwax8<���3%7|P��LnzI�kT��82�9!&���S+e#��]�r�t8� @V��	�4�ڟ����p��W�߉+��2�=��ݒ�w��nR>���b��&��� �ɽ�*<e���8w��k�cp�l���N.�b��q~1��ɽ�*<eR�n�@�O&X�aҥ��0ŻA�y\Z٩G,(�Ě��δ8?Cv��p�.�����������y�ճ��}�����;��F�t�e�dA������q~1��ɽ�*<e�VJUT���M�{�Z�1.�ez7��������(-�hm��>0<S����~�p����^�+�E�Vl�q���������S ��V�����y�ճ��ȩ�Ļ�(�z~�(� 4��JZe��1� �����Ŀ�O��gSy���a�}cm�&*�q���������S �L��<$&��-Dc�����^B%�y�c7,?-�Y�������bC�x���b��6�-4�)�_π|UT�����^B%4�@_t����Qݓ˟s4�)�_π ����������'�e������Ki��Z0B��#��J���p�����5[1.c�CǼ���#�����x�};�����6�.���,�.��W���Z0B��"�ĥ�@�p������R�	�	0�CǼ���#���RD�R};�����]���9����.��W�|�	R��-Lċ�LY-.fyp�5�o���v�81�++����
�6�c� ��Uٿ�ю��8���&���N k�I9^�ï�Lz�K�R�H�]�ͻlU�� <�ZBgT��@,j ��8۬ȴ��j�Tu?4��p���w�ae�Ӏ4�;�Q��}8�*���x�)�[����u���̹尮l;�j��ɽ�*<e�
v�ƒm�9(ύ��Bɽ�*<eɽ�*<e����n��rɽ�*<e^��
:�*�)��Y�*B������."1Do�zR�J}����q�����e��1� �����Ŀ�OñiE����nL���xr��<I}��,�����}nUD�DD#�˴��56��@�� ���q|���)u/��L�<Q�]�Q�MY[v�_�>[��H�����!�����V8ߊ{Hw��	�;�;�<�ɠ)�F�����+���G:fGv��l���SI�\U�>:�����n��rɽ�*<e���U�&4�K����!<�NO'�"�d�;�@�j/�j��ڭWH����	�;�;�M
����ɽ�*<e�����+�n�/�Gg��	� �Ei�OϿY�f�af�w��Y�3�9��F�t�e�7��r|�.�YС�VJUT���?�(<����vVK�`���;�	Ei�OϿY�^|��]`�Y�3�9��F�t�e�7��r|��v�1�V��VJUT���?�(<����vVK�`^|��]`��,����������Ղ5�7��dh��@�� ���q|�����rq��&�������Y[v�_�ɽ�*<eN�����K5�B���>���i3�^��P�6;7}7|P;���\���ֻ'i��\;�&��z�IYLy�h��ҝ[��R�ɽ�*<eD���p �W"!��ٜ;>���i3�^�Д�٪,=~�����\���ֻ'�ȡ�X0���b\	y`��h
�K=4ҝ[��R�ɽ�*<eVd������ʴCj��i��\;�&4�)�_π}��X0��j��Eh��)V���U`H��,4���?w���J�����FӖ�^(�C�@� g�+�����ʠ��6M�TqSݲ֕���w�u��Q�)y��Z0B���z&Ƙ�����#ڄg��1-P���h
�K=4ɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e���r�<,�����]��ƚ���b�	��*SD�G�9#Rz�g��Oa�׻\-�!���-l	*vY[v�_�ɽ�*<e7��� hE,>����$���h�%���N�-������K�P ��謋:M�TqSݲR1�#P,ޖ�,�\������ɽ�*<e8���pe��] �, �˞Q�Z�[4˛��O��]�� �??�8�|q{+��hM'��INd�N���ɽ�*<eɽ�*<e��]/߷�W�߷G�ey/�K�?V��{Y\iq�tQ��C�q�X�<QPmssU�*N6���^���T���V�!GA>>�-^wq0�Ks�b� �+�+o��[}[��z��I-��c���Amg�{��Uq f�&��q�"I!���P>�=Z�'[P�u�1? ��6�2��p�ɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<��ɽ�*<e-��fΡ��k��4t�p�(�Z��a��-�hm��>0s���Q���?�*���H�b��
L���y���C������ɽ�*<e���Dx�v�Or���Jv%:�Q_�E�\*
�-=�QO��]�� �??���	�d��@��M����0�1�ɽ�*<eɽ�*<e���b?Tw�\Jm�Q�8;7v����Ne�D��ܗ	�4�ڟ���
�(G�y��5���c�H�hoM�,K�%-
+[ɽ�*<eɽ�*<eD���p �WZ|[s%�o4q��t�kRIꐦO�j���}O���Nc�T���֤�T��U>��T�N������B�C�q�X�<Q����V
`�c�A$���ꈍHg�8�3�F��7u$�򝧭9l��ג$OJ�7�^	$,�_�����@�]�H۝���+�Jr����&6ɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e:j���+�oaf�	��,Jr��v@�0ܜ�����X�aҥ�����&g�vn���N.�b����Ǆ{� ̛#ɽ�*<e�i{ޝ��i�[.�[���3�Cz�^m��"�,w#Ne�D��ܗ	�4�ڟ���
�(G�Ɖ�D��0L\[5���d�NM{9q��ɽ�*<e�"�|��(��%�>v;��	f��Աl���#R�b����(O%��;!��;K�Raz��w$o��3b��ʼ�?�(<��ɽ�*<e!�T9�u�P�+H�"��i�5�kD���&�Kq��2V���,."�9A�F�m �
�HVH<������n��r���}O���Nc�T��w�~Ġ��`����T�t�=	E���;�V�
%�n�>�B"b��i���sX!䖸3���̹尮l;O��a[��=��X��cQ�]�Q�Mɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��ܑ��h"z<�'~�� _�5yo�Xꦻy~�q�����u���������p`�ժH���NM{9q��ɽ�*<e`ύ���#�, ��T�"#��K�d��C !b����(O%��;!�ٖ�3������%O���f��t��?�(<��ɽ�*<eD���7�7��;�d ��D���p �W3?h�������^B%C=֡��́��]-����P�6;7}Q�D�.�^ɽ�*<eɽ�*<e�����^�*C���w9:w��a]�x�r%=YF�u��}V�A�iz�'kL�9�6� ?�hy�}�/WB��,."�9A�F�m �
�X<Ҹ(ML��9q:Xx3���^���.�ř���WJ������]�ͻlU�Å�2�*���yot��;���ǋ'H)�@wV]��%�ɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<eɽ�*<e^��
:�*�~�sh-�߮� ��V��(�틪��W=.�A\����������#(�ZZZ���?�(<��ɽ�*<e����F�i���!`�ۄ�%�>v;�?�&�$�(���^B%C=֡��͡u�6�f�3���
���2�'8{ l��ɽ�*<eɽ�*<ejG�7�7�okx� oK��:�����
Y\�er"�꺯z^kM�m��X�s�Q^ڝ����%�:ҝ[��R�ɽ�*<e+�n�/�G/���?��?ň?���.:-|N���G2(�|�:霐��{ѧ���9HO��.�[���vR�HN^xΊ�A�iz�'k�At����i�0R#1���9a�н�r����ʻ�L �j\?����Q� ���Ɯ�h�Ī��G̐>B�n�����Xv�k��=!��(]��s�kɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�G�x9��FE�&I��}�, ��T�q�=� ���=��od9�ܳ���-V'Ba6j�sk��x�\�uɽ�*<e��_��l���<I}�^�u�G�f���l�@���
Y\�er"�꺯z^kM�m��qc'|*�}�o���ҝ[��R�ɽ�*<eNȾ5TDΔm��ڴg���;�V��#��3%7|P��LnzI�k�
T������8��n�:j��ɽ�*<eɽ�*<e���U�&4�K����!A*C�x&�yh�S
cP��yQ^sU��m�q&��a�]mZ*�->B^A+kK�ȹC:霐��{ѧ���9H`S��|��uZ1����k�I9^�y��a�Ξ7��ɇ�F�b=��K�X�j�^��$A9�+�RU� 0��%rw�;L�::^�Q��	�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�4����k���A�X:蕵��X�x�!�I�mek�cp�l�AѼ]'�~�!�*�X�I�� �pҝ[��R�ɽ�*<e�}��^�|"y�׫&�(�rv�����h�]l�3%7|P��LnzI�k�s7�}��/���>;�#k;���A��ɽ�*<eɽ�*<e��I��㱡 4���:o/���?��"��>�w�f��K�����H�گ�`�\�m0a�/���?��iE����nɽ�*<eɽ�*<e7[��İ��jN�̓���׀�.H���?��B��}X|W?+~I�)�]���y���/\��MPW��~h��c�6U��m�q&���^���$q^�.�2�9��z-����hԚԾ3��R
y�h�ᕑxpu��8B`}���$�y��k��dU'ѳ��w���
v�ƒm�9(ύ��Bɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<eɽ�*<e�MO�~Iy'p�k㐊��;0>(�z~�(� 4��JZe��1� �����Ŀ�O�1wg�i"yPɽ�*<evS+ё@�˴qZ5�+�/I��/w��\��"��>�w�f��K�����H�گ�` �D�O�h>)u/��L�<�K�{b�&ɽ�*<e�p\�Ì����z����xz��������������K�P ��謋:M�TqSݲ܎h*�Gm�v[o�I�^�����ɽ�*<e�H��g澚c����T0��e��g8j�R���	u|4���V�!GA>>�-^wq0�	⏌��n|����e½8����~I�)�]��wl�=P'�#^��׊� g�+�����ʠ��6�V�旾sb��i���sX!�Ɣ}Y��� 0��%rɽ�*<eg��1-P���h
�K=4ɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�G�x9��FE�&I��}�, ��T�<���^�jT(�z~�(� 4��JZe��1� �����Ŀ�O������?�(<��ɽ�*<e����F�i���!`�ۄ�%�>v;�?$�r�|�3%7|P��LnzI�k�F{N.J��@��M��|���n?�(<��ɽ�*<eD���7�7��;�d ����j��G$���-�6�b����(O%��;!�ٷ��{�}f�ϯ�㳔J�����?�(<��ɽ�*<eșQ�z�~��$�\׉���4ł���Y����zݝ3%7|P��LnzI�k�F{N.Jɥ]�gk~�/����?�(<��ɽ�*<eșQ�z�~���;=6
��u��_^A����6�aυ����K�P ��謋:�V�旾sA��y^G��B���b�ҝ[��R�ɽ�*<e+�n�/�G�_�av"c돦��v�5�'��,��"��>�w�f��K�����H�گ�`vP�����c�H�hoM�9�<7���ɽ�*<eɽ�*<e�����^���J�= ȉ~��?0��l�FD�V����B({C�q�X�<QPmssU�*N6���^����n��r���}O���Nc�T��w�~Ġ��`����T�t�=	E���;�V�
%���7�1�b��i���sX!���7�1�̹尮l;O��a[��=��X��cQ�]�Q�Mɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��ܑ��h"z<�'~�� _�5yo�Xꦻy~�q�����u���������p`�ժH���NM{9q��ɽ�*<e`ύ���#�, ��T�"#��K�d��C !b����(O%��;!����7�1����%O���f��t��?�(<��ɽ�*<eD���7�7��;�d ��D���p �W3?h�������^B%C=֡���A�O����忘P�6;7}Q�D�.�^ɽ�*<eɽ�*<e�����^�*C���w9:w��a]�O��'?�U��A�iz�'kL�9�6� ?�hy�}�/WB��,."�9A�F�m �
�X<Ҹ(ML��9q:Xx3���^���.�ř����:#�u]�ͻlU�Å�2�*�3����ue�;���ǋ'H)�@wV]��%�ɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<eɽ�*<e^��
:�*�~�sh-�߮� ��V��(�틪��W=.�A\����������#(�ZZZ���?�(<��ɽ�*<e����F�i���!`�ۄ�%�>v;�?�&�$�(���^B%C=֡���)�ߙmit����
���2�'8{ l��ɽ�*<eɽ�*<ejG�7�7�okx� oK��:�����
Y\�er"�꺯z^N�� �� �?��R���:�����%�:ҝ[��R�ɽ�*<e+�n�/�G/���?��?ň?���.:-|N��Wp 	�F
:霐��{ѧ���9HO��.�[���vR�HN^xΊ�A�iz�'k�At����i�0R#1���9a�н�r��������r��Ub��i���sX!�o%�;�bZ�'[P�u��/���%��X��cQ�]�Q�Mɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��ܑ��h"z<�'~�� _�5yoq�=� ���=��od9�ܳ���-V'Ba6j�sk��x�\�uɽ�*<e��_��l���<I}�^�u�G�f��-Ȳ�N�#"��>�w�f��K�����H�گ�`�ɜ��8���}�o���Y[v�_�ɽ�*<e�p\�Ì����z�I��;˽�񊅄NＡ_�6;�B��K�����H�گ�`oc�v^���"C�ӀNM{9q��ɽ�*<eɽ�*<e��j��G$8�2Z�Jt0#@}i�q�
Y\�er"�꺯z^V9��V:=�I�`�q���v�1�V�ҝ[��R�ɽ�*<e+�n�/�Gi���!�)��'�9�<��;�sNe�D��ܗ	�4�ڟ��]��Maz�����RP��;J��>,K�%-
+[ɽ�*<eɽ�*<e���d����ؔ�����8;7v����?�&�$�(���^B%C=֡����=H��A��c�H�hoM�9�<7���ɽ�*<eɽ�*<e�����^���J�= ȉ~��?0��+�
�n�ޱ�C��QA�iz�'kL�9�6� ?�hykK�ȹC:霐��{ѧ���9H`S��|��uZ1����k�I9^�ï�Lz�����K�P ��謋:b��i���sX!��
Y\�er"�꺯z^�z&Ƙ��=�Y�����#ڄɽ�*<eɽ�*<eɽ�*<eǋ'H)�@wV]��%�ɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<��ɽ�*<eɽ�*<eɽ�*<e�KzM|��,������<�X���K�o��c�hz�;3��PY���F��
�W���[�&U�,�5�(�z~�(� 4��JZe��1� �����Ŀ�O��h
�K=4����kc靯�;�4�)�_π ����������'�e�j|�2�F+f���kY�`χ�a$����^�M�"�ds��R��6G�2�K�����]vm�r�7�k�cp�l�AѼ]'�~�!�*�X�I�� �pY[v�_���7�1��W���[�&�E�?9D�uǎqh��˴qZ5ت�$��NCZ��F�t�e�c���L)�/(T�F(��ɽ�*<eɽ�*<e�����+���G:fGv�ݹE�=5�4QOB-�y�ɽ�*<e,4���?wɽ�*<eɽ�*<eɽ�*<e�� �3Y�S���ʊH�Δm���7�U|�V�ΗCf�|���R���7��$`љR�ɽ�*<eɽ�*<e�������i�OϿY�M�L>�;>cc��R��Mbɽ�*<eY[v�_�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��{P���� <�t-*��,������G:fGv������6�\� R�E��ɽ�*<eɽ�*<e��@�� ���q|������g�#wF��@�OG�ɽ�*<ex�\�uɽ�*<eɽ�*<eɽ�*<eɽ�*<eY�I����b\	y`��,������G:fGv�C�b�MPɽ�*<eɽ�*<eɽ�*<e��@�� ���q|���0ڧ�AO4ɽ�*<eɽ�*<ex�\�uɽ�*<eɽ�*<eɽ�*<eɽ�*<e!�T9�1����X���F�t�e�'l�����d�!I�2ɽ�*<eɽ�*<e�����+���G:fGv��l���SI�\U�>:�ɽ�*<e,4���?wɽ�*<eɽ�*<eɽ�*<eɽ�*<e+�n�/�G/���?���,������G:fGv��l���SI����!�ɽ�*<eɽ�*<e��@�� ���q|���/���?���AE
!�ɽ�*<ex�\�uɽ�*<eɽ�*<eɽ�*<eɽ�*<e!�T9���z�IYLy�oc?3�<ڭWH��;��)����'d����ɽ�*<eɽ�*<e�&�JG��b�j��EhV�v�Ee��h
�K=4ɽ�*<e�VJUT���?�(<��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����I>���i3�^���q|���i���!�)�49�iv (ɽ�*<e�/���%�\���ֻ'^{�1u$�J_���Q�]�Q�Mɽ�*<eNM{9q��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��r���
�JP$��k3�:R1�#P,š�	"�$ɽ�*<eɽ�*<e@�j/�j�������K�P ��謋:M�TqSݲR1�#P,ޖ�,�\�ҝ[��R�ɽ�*<eɽ�*<e�W7P�%7��ɇ�F�jG�7�7��!�/f�O�8�|q{+��hM'��IN�������ɽ�*<eɽ�*<e�a��aO��]�� �??�8�|q{+��hM'��IN�v�r��?�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e+�n�/�G/���?��Qq�t��V�����=�w��\��ɽ�*<eɽ�*<eɽ�*<e"��>�w�f��K�����H�گ�`�����=�)u/��L�<9�<7���ɽ�*<eɽ�*<eɽ�*<e�@���������ݣ�;�d ���k3�:��e��1
�<�ɠ)�Fɽ�*<eɽ�*<e@�j/�j�������K�P ��謋:M�TqSݲ��e��1
��v[o�I�^ҝ[��R�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����^��Q/���t���̌/���>;�##�˴��56ɽ�*<eɽ�*<e?$�r�|�3%7|P��LnzI�kt���̌/���>;�#��g���?�(<��ɽ�*<eɽ�*<e1稆���%��+ v����%�>v;�Qq�t��Vڇ��C�/���?��ɽ�*<eɽ�*<eɽ�*<e"��>�w�f��K�����H�گ�`ڇ��C�/���?���'8{ l��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e!�T9�u�P�+H�"U'w{cy�eAΣi0���-Ȳ�N�#ɽ�*<eɽ�*<e�/���%��
Y\�er"�꺯z^kM�m��AΣi0���}�o���NM{9q��ɽ�*<eɽ�*<eɽ�*<e��3�����|t����A|���ϝO�}���8���b��M&ɽ�*<eɽ�*<e?$�r�|�3%7|P��LnzI�k�ϝO�}���8��/����?�(<��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eD���p �WGӛ��x�5�u�6�f�3���
���2ɽ�*<eɽ�*<eɽ�*<e?�&�$�(���^B%C=֡��͡u�6�f�3���
���2�7F'�]hɽ�*<eɽ�*<eɽ�*<exP�Z�W�SF�W��A��] �, U'w{cy�e�X�s�Q^�5�'��,��ɽ�*<eɽ�*<e�/���%��
Y\�er"�꺯z^kM�m��X�s�Q^ڝ����%�:NM{9q��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��]/߷�W�߷G�ey�/�ӄi�4���%O��(T�F(��ɽ�*<eɽ�*<e���E�֦$b����(O%��;!���/�ӄi�4���%O��'~_�~N�����ɽ�*<eɽ�*<eЖ��ٿEe���I���z��4�l	}�I�b�H濘P�6;7}49�iv (ɽ�*<eɽ�*<e?�&�$�(���^B%C=֡���I�b�H濘P�6;7}�3\�]P�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�H��g澚c����ٹB��ZY�r)1�ڹ�m��"�,w#ɽ�*<eɽ�*<eɽ�*<eNe�D��ܗ	�4�ڟ���
�(G�r)1�ڹ�\[5���d�Y[v�_�ɽ�*<eɽ�*<eɽ�*<e��Z0B����%h���� 4���:o��?��Bⴹ�w$o���!I�2ɽ�*<eɽ�*<e���E�֦$b����(O%��;!����?��Bⴹ�w$o��w�	�6�c�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<e7[��İ��w�f��=�m��3+� ���@��M���>Է4ɽ�*<eɽ�*<e�a��aO��]�� �??�m��3+� ���@��M�zA�Lɽ�*<eɽ�*<eɽ�*<e�2��9�|nE�d��OhΔm���ٹB��ZYΫ~u��18;7v����ɽ�*<eɽ�*<eɽ�*<eNe�D��ܗ	�4�ڟ���
�(G�~u��1c�H�hoM�K�{b�&ɽ�*<eɽ�*<eɽ�*<eɽ�*<e���U�&4�K����!���I����%O��(T�F(��ɽ�*<eɽ�*<e@�j/�j�������K�P ��謋:�V�旾s���%O��'~_�~Nҝ[��R�ɽ�*<eɽ�*<eɽ�*<e���{�}fjG�7�7��!�/f�O�-KB�i�&�ӂ[uɽ�*<eɽ�*<eɽ�*<e�a��aO��]�� �??�-KB�i�"���y��,4���?wɽ�*<eɽ�*<eɽ�*<eɽ�*<e+�n�/�Gl� �J�ࠓ�I���w$o���!I�2ɽ�*<eɽ�*<e@�j/�j�������K�P ��謋:�V�旾s��w$o��w�	�6�cҝ[��R�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����^��Q/����F{N.Jɥ]�gk~��b��M&ɽ�*<eɽ�*<e?$�r�|�3%7|P��LnzI�k�F{N.Jɥ]�gk~�/����?�(<��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�4ł���w�f��=�-KB�i��
��nE�y;�<�9�ɽ�*<eɽ�*<e�a��aO��]�� �??�-KB�i��
��nE]C��u<ɽ�*<eɽ�*<eɽ�*<eɽ�*<e+�n�/�G�_�av";�h��}��N��@��M���>Է4ɽ�*<eɽ�*<e�a��aO��]�� �??���}��N��@��M�zA�Lɽ�*<eɽ�*<eɽ�*<e�2��9�|�Tf�^eVΔm���+f���kYK��Ak�28;7v����ɽ�*<eɽ�*<eɽ�*<eNe�D��ܗ	�4�ڟ���L�KJK��Ak�2c�H�hoM�K�{b�&ɽ�*<eɽ�*<eɽ�*<eɽ�*<e���U�&4�K����!�:�;�n�T̨̻v��š�	"�$ɽ�*<eɽ�*<e@�j/�j�������K�P ��謋:��9�E"McT̨̻v��ޖ�,�\�ҝ[��R�ɽ�*<eɽ�*<e�W7P�%�����x�jG�7�7��!�/f�O�
j����hM'��IN�������ɽ�*<eɽ�*<e�a��aO��]�� �??�
j����hM'��IN�v�r��?�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e+�n�/�G/���?��Qq�t��V�ɜ��8���-Ȳ�N�#ɽ�*<eɽ�*<eɽ�*<e"��>�w�f��K�����H�گ�`�ɜ��8���}�o���x�\�uɽ�*<eɽ�*<eɽ�*<e�2��9�|�S<��伸��;�d ��eA�-�\ձ�ϯ�㳔Jɽ�*<eɽ�*<eɽ�*<e@�j/�j�������K�P ��謋:�x�A-���ϯ�㳔J�h
�K=4ҝ[��R�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�]ӞvQq�t��V�	�
�W�5�'��,��ɽ�*<eɽ�*<eɽ�*<e"��>�w�f��K�����H�گ�`�	�
�W������%�:x�\�uɽ�*<eɽ�*<eɽ�*<eɽ�*<e!�T9�u�P�+H�"����p.�I�`�q���|�/��=1ɽ�*<eɽ�*<e�/���%��
Y\�er"�꺯z^V9��V:=�I�`�q���v�1�V�NM{9q��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��r���
�JP$�eA�-�\ձ��Aau�]��H�Q�Bɽ�*<eɽ�*<e@�j/�j�������K�P ��謋:�x�A-����Aau���9�eSpҝ[��R�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�e��\ȟ�:6H�� ����&�5tXCB?�<X�aҥ���4f<W��ג$OJ�7��D����H��
�����1����bT�>^Gʵ���2�#h�)�r���PY����*�U�2��T�\�To�ǭ�4%Γ�?�I;�68�Fxɽ�*<e�i��K��������zU?��4�Yz`E]��~)��Θ[{����vL�)������U�8AmI�z�#-K}���5�l#�ѝ�j0t&r��/?���hh�ro���İ�A��SƁ�7w�'m�K=�_��2G:����)�Lw��g']5��kL���RI?�fm%�Ef�9L��P�a��D��VZF��m��N�N�W\�ߐuX�q�����V��U?��4��<�����.���)V�T(�<7���_P!_0��X^��U��h���Lw��g']5��kL���RI?��A�b��3L��P�a��D��VZF��m���&XOD��ߐuX�q�����V��U?��4��Fzΐb�.���)V�T(�<7���_P!_�BC�S�U��h���Lw��g']5��kL���RI?ά�BM��qL��P�a��D��VZF��m��/��$"���ߐuX�q�����V��U?��4���W��\Ź�.���)V�T(�<7���_P!_�hb�B�_ðU��h���Lw��g']5��kL���RI?�����OAL��P�a��D��VZF��m���'4�%�bD�ߐuX�q�����V��U?��4�K��k�.���)V�T(�<7���_P!_�a`�;��U��h���m �"}�r���PY�֏��-��)ӕy��-�+�F�X�aҥ���p�#
�!�<�DR��#NgG�g'ë�Ꚗ��1AiDQ�]�Q�Mɽ�*<eX���Ѯzꏼ�t�_��%�6��fAϟ�o�	� ����g\���ֻ'i��\;�&4�)�_π�m����톣Z���-\d*C�S*���/��`����#ڄa�磅"��Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<e�����^��
:�*�~�sh-��:\��lRˋ_�^l8>s�=��od��)V��H�b��
L�^0�\<ef���N.�b�j|�2�Fy'p�k��0n� �¾^1�?q�-ɽ�*<eɽ�*<eɽ�*<ej	�%w\�����mq[0�<�(p�>u�b�Px���P��MK�s�Zɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�fy'p�k�.	o�L��S�;��$�Q�]�Q�Mɽ�*<eɽ�*<ej	�%w\�����mq[0�<�(����s��^�+ �0��MK�s�Zɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�fy'p�k�ϔZ��S�;��$�Q�]�Q�Mɽ�*<eɽ�*<ej	�%w\�����mq[0�<�(�r��m� ��+ �0��MK�s�Zɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�fy'p�k�v��[��S�;��$�Q�]�Q�Mɽ�*<eɽ�*<ej	�%w\�����mq[0�<�(V��k��̖+ �0��MK�s�Zɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�fy'p�k�T�fe;�QS�;��$�Q�]�Q�Mɽ�*<eɽ�*<ej	�%w\�����mq[0�<�(�_(L��c�+ �0��MK�s�Zɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�fy'p�k�B�a\1	nBS�;��$�Q�]�Q�Mɽ�*<eɽ�*<ej	�%w\�����mq[0�<�(���?+�@�+ �0��MK�s�Zɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�fy'p�k㣚m�Y���S�;��$�Q�]�Q�Mɽ�*<eɽ�*<ej	�%w\�����mq[0�<�(��j0��;�+ �0��MK�s�Zɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�fy'p�k�=�f?u{�S�;��$�Q�]�Q�Mɽ�*<eɽ�*<ej	�%w\�����mq[0�<�(#ɀ}�&>i�+ �0��MK�s�Zɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�fy'p�k��ϴ�@�S�;��$�Q�]�Q�Mɽ�*<eɽ�*<ej	�%w\�����mq[0�<�(py@2a��i�+ �0��MK�s�Zɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�fy'p�k�pF�3�[9~S�;��$�Q�]�Q�Mɽ�*<eɽ�*<ej	�%w\�����mq[0�<�(p����^��!�Tn�PMK�s�Zɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�fy'p�k�.	o�L��71OyƧ�<Q�]�Q�Mɽ�*<eɽ�*<ej	�%w\�����mq[0�<�(p����^��9	k�ⴆMK�s�Zɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�fy'p�k�.	o�L�ߞAȢ��6Q�]�Q�Mɽ�*<eɽ�*<ej	�%w\�����mq[0�<�(p����^�?��f�,݇MK�s�Zɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�fy'p�k�.	o�L��Q'f�<�ZQ�]�Q�Mɽ�*<eɽ�*<ej	�%w\�����mq[0�<�(p����^�*p_	�R��MK�s�Zɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�fy'p�k�.	o�L��:�B��&�Q�]�Q�Mɽ�*<eɽ�*<ej	�%w\�����mq[0�<�(p����^�\��Y"~�?MK�s�Zɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�fy'p�k�.	o�L��X!���5IEQ�]�Q�Mɽ�*<eɽ�*<ej	�%w\�����mq[0�<�(p����^�;��8G(MK�s�Zɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�fy'p�k�.	o�L���9��3(�ɽ�*<eɽ�*<eɽ�*<ej	�%w\�����R
�CI���$�$�w�'� �۟�6 �D�G�9#|�����N���Q�)y��$�-�bJ	��$�1�x0Ycɽ�*<e���[��<��;τ��2������7a~�	��1�z�'G�7�߰XnVC4[!7,���f���xɽ�*<e�:�<�.�ؗ���v��_P!_��~��7�q�Xm.��ߐuX�q�g']5��kLDQǺ��@y~�^+���B�j�^9/-E��+lJ@Ҷ#�hMU)�_>%"	�E׋������z�{Ά�[����;(�Y�>���?�L��P�a��D��VZF��m���|(~��
��ߐuX�q�����V��U?��4���[���A�.���)V�T(�<7���_P!_h�Ү����U��h���Lw��g']5��kL���RI?��U���v�L��P�a��D��VZF��m��-��y�����ߐuX�q�����V��U?��4�J�����.���)V�T(�<7���_P!_�6�̚r��U��h���Lw��g']5��kL���RI?��g�.@L��P�a��D��VZF��m���LD��@�ߐuX�q�����V��U?��4�H���.��.���)V�T(�<7���_P!_��6��kP��U��h���Lw��g']5��kL���RI?�����X0�L��P�a��D��VZF��m��V�D�����ߐuX�q�����V��U?��4�sXi��L�F�.���)V�T(�<7���_P!_̅�k=�g�U��h���Lw��g']5��kL���RI?�)nV�i�(�fkN�F��&B�B_E�U?��4�*��@M�aU{� P����(�틪��W=.�A\��5�r�鐦D�4�i�K�ؽ->*W�����Mp冚aɽ�*<eɽ�*<erL۪w�Ib�D�4�i�K{��%B{$Jr��v@�0���Wnh����@�� ���q|��������I�� �p�VJUT���U���N�*�o]��_��*�ɽ�*<eǋ'H)�@wV]��%�ɽ�*<eɽ�*<eɽ�*<eNM{9q���4����k���A�X:�!]�?T�R���~�I(�z~�(� 4��JZe��1� �����Ŀ�O�����S��i!���H9�����Pwma=� >*��������l�ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곬��Pwma=ѷ��G��-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곬��Pwma=���w̜�-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곁<�DR��}�+�IO-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곬��Pwma=��1zs9�-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곁<�DR�~�<����e-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곬��Pwma=����w%�-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곁<�DR��N�{3E-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곬��Pwma=ڀ��C	�-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곁<�DR���)�)5�-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곬��Pwma=aj�H����-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곁<�DR��`?�ƶ�-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곬��Pwma=��aC`-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곁<�DR�>�g۴p�-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곬��Pwma=���q�]�-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곁<�DR�Ǎj��c�-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곬��Pwma={ZN �w-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곁<�DR����p=ߞy-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곬��Pwma='��3��NG-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곁<�DR����BF�4�-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곬��Pwma=ex�
�Mn-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곁<�DR���W�r�#"-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곬��Pwma=�j�+���-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곁<�DR�}=���/�-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곬��Pwma=�.�It[�e-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곁<�DR�g�����#-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곬��Pwma=Ԝ��a�-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곁<�DR�ɲ����-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곬��Pwma=6�6.Hb�#-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곁<�DR�q�,��R-&J�� ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곬��Pwma=Cᮦ�ɤ�K��c��ɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wY�@o��W��-P�ġ|wu6��Zl�e`Wb֢�<�����e���w�\
h�["M6f��������5�JF�M�Vy�cgͼ��UQ�N��V��G���Y���C��&�-�,�X�Ÿ�f�2_B@:P��dS	nT��e�&��F]�J�������	U�֝�%��LP�b�I�hS\'��/���`b]P�L��ϰ�9_��]-͍)�,\���� I���X�%���=��dn'y&̢���N���ꗳ�)�70bxN7~/Ǧ��!Fȵa�E�UJ̘�P���W��-�\��\����WgƘc���Jt���M���bf�\c�ꗳ�)�7�;⑤���a,�"�빱x�Q<�^eg��ɂ����c_�o� x/���C $P��!zsv|MC�[��ĺ6
&���?��������Y���i{\�M�Q#�`>�P����Yy��0�	ĭ��n�W���\?�R�?3�h0)�E�Z��(w
�7`�	�6'�����<5���K�����,%GJ�k���.Ҋ[m]1��F�^v�'-Ɨ�8;�gi��{�]<�S#��B����2"��
��V������+�v��Tj0��L�m��7���dO��H�\?�4x!�i輸m�a��&�^��=3���,je6�����B�g��o&76� ���+ɾJ�Y�WX���v�	p��i���y�6]v��P|Λ#�2�[�k�tf�����0U������J�yP��}H�{_�.�@)1�7-��H�&��_�6�*�q#�L
2�������̹�"�j��;�kԐH`�Q��
I�DYZX�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��?h�Z����Up	ȶ5�|d$o����5�l�ɜ� 1"�Op�ű�!� Sv�0.���&D�HF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8����T%�g')l`�AG�0����9�)�Txi�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8���W�|�Z�p���	j�֏�"%��e.i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�@�ae�� >A�Pɔ=Y3���ڎX"����ݸ8؋ֵ|�����N���Q�)y�o+�����Uj+����1�2P'L���Ę�c(W'4�l&ꬶ�R�G�x9��F�G��/�gj�X��]��zN�����ɽ�*<e�.��W�Hv@�����Uj+����}NВີ��/�žC����N�������Zƚ�������]��5�F��7 Z��I�D�J�ɽ�*<e�x[���K&��06(���� ��#*sīX�(��O��xx�yN�F�8I5��Oh`B�VT�́ɽ�*<e�(���V8��+ Z���cW� �ϵ%[��zN�����d*�cHа���<���^.�+:-nPC"Ɔ�;��t�^	�ER���-��Ę�cw�)3��Z��������3�jh��kE�ML�ic��ݤ���S���)�ɽ�*<e91��?����06(�����N���sīX�(���I�e�H�KV��iI]�P�.�F{T�_0���ɽ�*<e�g?k�Vtև̸B����NI|	*���W<:KRKD�vQF���&B���V��P ����X���}�,4���?wʉ$�Hl�/�%�M!O��y�2f!����N����j7�po�1o�Z����\�?�5��Oh`B�VT�́����C��/���?�䕢�cW΁��Җ LF�zN�������ky�-�땢�cW΁��Җ LF�zN�����0�����ʨf��w<����N���3��͠��1 K��0�||�,�h{���{ z_.?�P!����Si�M��GW�yN�F�8I5��Oh`B�VT�́ɽ�*<e��rq��&(�xt��:[�yl2����ar��Z�.vS+ё@�_d�Ǹ����<�i}�E��7ۅ��v
ZF�N����4���/���?��N�
�I���Z�������r�_`�m���dv����A)�^U�ɽ�*<e���p�S?��h�Ki����|*L���,���w��d���������A)�^U�ɽ�*<e0�J����6��U��RKD�vQFO@�����w��d��#��k�2u�>��d�F��[�I�T�i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S�A�b��d�1�p~rևl�4��wy f��F=�����F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��5�� �(д�`8�1�ڹQM7HW��MyޡP�3<N��lCƵ%��hb;��8�*���xbIF�L3R��N���CƵ%��hb;��ۭY��'�K-���j̧th����CƵ%��hb;���&�=��ɽ�*<e��~^-C�tPfW��Xƻ�2��gƧ)������M6��M�0���=x���]L�Eɽ�*<e��#��HP8����մ�ob��i���sX!�nZ�9��Iɽ�*<e�ҋ\�d����#ڄɽ�*<eջY@f����cW�ɽ�*<e���˺�1�}U������/���%󬖃�1AiD���cW�ɽ�*<ea��%�IO��:��*��/���%�F�W���ʃ��V�uCMɽ�*<eR㠍�������-�ɽ�*<e�T�=fR{��+�Cp6ɽ�*<e���`����!I�2ɽ�*<e�� �QȦk�v��ɽ�*<e���`��������d<������of�z�ΙA�̸B�����{���̙ɽ�*<e_�@2z���"vЅ\��a�k|jZ��˪��D�K�am@�G���L�w�ɽ�*<e:���)�9�š�	"�$ɽ�*<e`4BFB1T��y��ݓ�ɽ�*<e���U�&4�<�ɠ)�Fɽ�*<eׂƯ78��QC��i���ɽ�*<e!�T9�"�l��Z=�ɽ�*<e�g׆������cW�ɽ�*<e�]Ӟvɽ�*<e�/���%�@0r���9ɽ�*<eɽ�*<eVd�����<Y��+�2����(��b\	y`����V�uCMɽ�*<e��r���|�/��=1ɽ�*<e[�!��QC��i���ɽ�*<eZi��LύE��9���wo�	h�[q��V��2��Aqz����p��ɽ�*<e7[��İ������!�"�Y�n���_d�Ǹ��݁W/���ɽ�*<e+�n�/�G5���.���i`X�F���~l�������ꖞ8���í�2ɽ�*<e�i75�����w��d�&ꬶ�RU����"���y������p��ɽ�*<e;^(���Ov�H��<\� <�t-*��@K��:�{v�H��<\� <�t-*�ھi��͗
��I�v�:����p���)�w׽�ɽ�*<e��nE�$,^q�O'z��b��i���sX!�A�=G�BHɽ�*<e�ҋ\�d����#ڄɽ�*<eջY@f����cW�ɽ�*<e���˺�1�}U������/���%󬖃�1AiD���cW�ɽ�*<e�#����Ǐd��-QJ�/���%�Awo��o�B��@ȏӽɽ�*<eg3�GIJ����P�ɽ�*<e+�>���4��d�B�:Yɽ�*<eUp"C�U �f��S�Hɽ�*<eU��p�>
zDS&63��ɽ�*<e+�n�/�G{M�y0��bm�B���6�:��D�7"�#F��8����T�����p��ɽ�*<e��.�΁���K�am@�؁)�yhڑG������r����T�����p��ɽ�*<eBv̾LB8;7v��������&B�Z�Y���DS&63��ɽ�*<e+�n�/�G*��F���Nd"�O����~l���ԏ0�i׈����p��ɽ�*<e�%(:�*Φ�-C��z����&5�w�������̵oc^~M3Y����A�Y��gc�0�I7�ɽ�*<e�8z�z@^�CC���q f�&�����������p��ɽ�*<e5���]�H������ꡜ��|�J���ϲ\�I72ɽ�*<e�}^B�Ņ�2O+�r�^�zsGN���o��
D�ɽ�*<e��Ҝ��������p��ɽ�*<e�ܧ��!�DhY��F�ɽ�*<eɽ�*<eջY@f����cW�ɽ�*<e���˺�1�}U�����ɽ�*<eɽ�*<eS�m}��W`��A��ɽ�*<e+�n�/�G�se]��T�R��RP^�ܰ��i`X�F��@K��:�{^|��]`�*�q�f��<ɽ�*<e�ݼY�ß��p�N5�E��<)�a�8�����/���%�5���.���S�w��Rd�ל
ϙ� ɽ�*<e�� ��V��n2���/^��"������R���7n=��>r��_ID�����R���7qu��8!ɽ�*<e+�n�/�G�se]��.)����p�qA��=	o�!I�2D{�S��c�H�hoM�a_ˌ�\ɽ�*<e��Z��d�!��Z�"٧[��C�IPd��Q����&B�Z�Y����h
�K=4����p��ɽ�*<e�������9���z�4�qt�M��Ϛ�9���r)"[
JΕO���ɽ�*<ej&W`�)�u:׈S�y��L��Ԝ�x���]L�Eɽ�*<e"����ݸ8؋ֵ|�����N���Q�)yzڨ�w���ɽ�*<e+�n�/�G���Xv�kɽ�*<eǋ'H)�@w���V�uCMɽ�*<eU��`���5��e�[v-%ɽ�*<e�p��V�e���V�uCMɽ�*<e���#�N�d��-QJɽ�*<e�^k��^[
B��@ȏӽɽ�*<e���`���..+`��ɽ�*<ewш�� ��3D>�d�ɽ�*<e_�@2z��Y��# N��ɽ�*<eZ:�?)HQC��i���ɽ�*<e_�@2z��"�#F��8#��U��Z6�Xz�T��!�(I����9�+�ɽ�*<e =s���GJ��tL:W������of��a�@��t���<���^��{���̙ɽ�*<e��m�����-Ȳ�N�#ɽ�*<el�жO$�5�;U��,1ɽ�*<e!�T9�5�'��,��ɽ�*<eC6�^`��8���í�2ɽ�*<e�H��g��Gܟ�ê.ɽ�*<eUu���B����V�uCMɽ�*<e��r��&ꬶ�Rɽ�*<ec�"�	M;�����p��ɽ�*<e)_�6-�p�\� R�E��/��JZ�+�W��#T���ڛ�*�ɽ�*<em�}����i`X�F�ɽ�*<e��e.���D8���í�2ɽ�*<e��vVK�`M�L>�;>cW1	tqtV~�nG�Eg2����㕢�cW�ɽ�*<e�����^�b2�M/��J�/���%�/���?��*�a���ɽ�*<eɽ�*<e�=X�Soj&��1��Фơ��� 3�^�&�����cW�ɽ�*<eՎF�)\k����-��/���%�91��?����+�Cp6ɽ�*<eg3�GIJY��# N��ɽ�*<e~�䓯���QC��i���ɽ�*<e�l�u+��v�ym��Aٰ���˫��J��=e��G5�td'3.�K(���ɽ�*<e+�n�/�GtseQ,�ٰ���˫��*ˋ���"vЅ\�.\~k:��zɽ�*<e�Xr��P�7ٝGy��;��f�vx&�@��A��mt�[Q>���ě��#��HP8����մ�ob��i���sX!���9%���kF�������2w��YE����� ��#*ɽ�*<e�:�#;��Ę�c5����_k`ɽ�*<eR��z��#�]� ��)!kF������!ڱ���sr��J�Zʛ5��M���>���6���&�|�D��x����Q���&�|�D��.�^<�
:�ɽ�*<e�x[���K&��06(���� ��#*�G�@9��ܻ�r�i:Mȅ�J�_��yl2���ɽ�*<e�&�|�D��"�#F��87U*���g�&�|�D��.�^<�
:�ɽ�*<e��X�ޒ-��F����ߔG�=��I��&6=��!4��Y5���&���W��5��M����Ve���\ꀪ�  �s郝��ɤF��7 Z��B�a�hꇲ��C��/���?�䕢�cW��Kn�:Ou
����.M-:���r���{72L%hQQ��p��u��d^��]����{72L%hQQ�wF�=d�Z!6��D2�P�����\�ic��ݤ����l�*�n|���=�^|��]`앢�cW�\�I;���ɽ�*<e��K�I4?�S��O�&�|�D��.�^<�
:�ɽ�*<e3\�!ќ�q�cW���c�0�I7�����n��r�7�'�\��M`t���<,4���?w~�V[��5T�e$̕T�:J�7�Bx��H!�b:eӪJ֐�f �a[����x�WoH0��T�d��2^���{72L%hQQ�s�������4���i���!�)ۂ%#B����N���6����=��8z�z@E�4k�G���F��7 Z���S���)�O@�����w��d��#��k�2��X��<�VC}�/��cF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^$��%�ㄕ�yд�";ν�BM��C��nhF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^nr�������w��U)��\��� �	Q�5�H"���b`�=c@�LT��~��!i��}�z�yf��r4����b�iؓ�"�JYw�8�r�rz����&��ל�y��}�!|�\X����{���Zݪ+i0�ɞ(�%��d�s�+��b7A�:�-��'�L����YT�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^Gm�I�	7�NC�Os��3Zʮml!c*�l�VUQ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��&Ic�E�,(r�p�V	�UVb�B��g��#E�,(r�p�V	 -ܒ�v�/���1b7N�ʆQ'�8���� ��E�5���L_ʻ�{�;D
'��`��b���<��'8��H��v���?v:@f�R�]��8z˷�����:�qڒ#-Դ���B|��;��N�ʆQ'�l�mf�E$j�P�@k)���T�M�V��4ud��E�p��u��dwRۣB����|}J®N�ʆQ'�ɽ�*<e�H��|��_�9I��>�װ�|�B� �aM�ZH�W��<Ƕ|���X�3{U5>g��u���B?O榼W��#T�{��8�L'6jE�،����)w����Zݪ+i�3H�����ɽ�*<e�~��gHQ�z =��ɽ�*<e"�s\:[YyA�fВ9��N^�P#�M�r?#���Aɽ�*<es����B8���C��=�?�",�ur�ӳ1�����ɽ�*<e�p�{��J�g�1A�)�������o:�]�ɽ�*<e�ԕOx�a,��?tr���4GH��͕A�������p��S�\�(�|�C:�����*����ܮm*���cW�ɽ�*<e��sH�L44Q�_nBY���D�-�7�C�!#% ɽ�*<e��oj�L���q��̿ ʅz�)Mͭ&<nr�m�ɽ�*<e��~�����O����P�����z =��ɽ�*<e��n
�/��*��E��UN^�P#�M�|!�K|�Vɽ�*<e4��؏�����]�!?�",�ur�����.��cɽ�*<e����[��"DП��S�łDV��޳6
Jɽ�*<e��ڈvV>�o�Zus|q�S�d蕴}3��3�	-����p�����A!q���"'�����*�� nx�6����cW�ɽ�*<e��O����k
UPֿ�u',�7�C�!#% ɽ�*<e����]�M/�Y.�P��|T�Xc���6�Ѻs�i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S�lR����鳫�Ț��5hEHX�����F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�W�	��g��e�F�Jx�r4'�qd!p*�~���M�,W)����z�"Uy��\=�B��YX��Ę�cd!p*�~�������,biISD�m��7���1�A��Ȯo�z�'4M���//�%
q�sڝ�o� }�DLc�w��6]�9������L����Ę�cr�����cδ�C:Z���/�žC����@��<�'!}��d��w����G��Mc__xZ��C�ɽ�*<e5���.���i`X�F��!TL�MUt���y�Pɽ�*<e0�J���QWk�HZ�s��l�s��\!����ɽ�*<e{R"&(ˣə�����x��F!��@z�Jɽ�*<e(z�E%x �ɽ�*<evE{��l��^5)��ɽ�*<e0�����&ꬶ�Rɽ�*<eM�3pI^C�����p��֪��"�+��bhF_ɽ�*<e�`F����A�Y��g�����>B�$Dɽ�*<eڜ�O�����NSad��kwO�&뿃m��"�,w#ɽ�*<e��/���_xZ��C�ɽ�*<e���L�8jɽ�*<e�!TL�MUt���y�Pɽ�*<eu-�!�J�ɽ�*<es��l�s����|��ɽ�*<e��u<@B�*G���}��x��F!��@z�Jɽ�*<eG�Y)S+�*G���}vE{��l��^5)��ɽ�*<e^��
�h&ꬶ�Rɽ�*<e�ܷД������p��f>>_YRcy�q<r�o�s&ꬶ�R�`F����A�Y��g�i{ޝ��i#-Դ�����p��ڜ�O�����NSad�����F+������Д�٪,����#�_xZ��C�ɽ�*<eXǿPÔ����	�E�X�!TL�MUt���y�Pɽ�*<ej�P�@k)���T�M�V�+D_/�����|��T��%zؕ��g�q\��/�žCkwO�&뿃���ft	������B!��Y�N:����p��ƚ�������H��8�M�3pI^C�����p���)�w׽�ɽ�*<e-H�x�k��В(��/���c�Ը��rJ�_C���>:䱠.�[bV��5F��4��A�Y��g�ŕI�(^�F��Ư@��=�5K�P�º>_�Ǣ��B?O榼W��#T��년�a�Ce���r�ɽ�*<eSE⫄ 2}
�E��d�4��R�ǹ��rJ�_C���>:䱠.�[bV�9P�Ɣ���A�Y��g�ŕI�(^�F��Ư@��=�5K��	܁hՏ���B?O榼W��#T��년�a�C�Zl��?_ɽ�*<e���+��C'�	�܉Jɽ�*<e��ڈvV>��jhD�TNk���,(nɽ�*<e����@��<�'!}��d��w���^�$��	t���l���rq��&�k0���ɽ�*<eɽ�*<e5���.���'d���������Ro��NSad��ɽ�*<e�+�r��y�ɽ�*<e"�s\:[Yy�v)���r�x���]L�Eɽ�*<eɽ�*<e�F�W�����#�t�X������Ro�C
�V[�ɽ�*<e�]�~���b\	y`�ɽ�*<e�ܷД������p��ɽ�*<e��}Gδ�-�o�c
����d�����#^�	�Nh��^Xɽ�*<e�
�9����ɽ�*<e�p�{��J�r�s��Ι��`V�f�Bɽ�*<eɽ�*<e��q�Ӭ=�u��OY�I#�L��~0H��r�dZɽ�*<eɽ�*<e;�>�"�!��Zb�Vq�e��d��m�� P�Hɽ�*<eɽ�*<e�\$�ǭ��;�3`-�$�:���f�G�6	6�Ƭm���r��
�Aɽ�*<eɽ�*<e���5$�bȇ�p��].й��|Ve\�L~�������p��'$��R��e�_o��u��ɽ�*<e�f�D ��dR��o-�}�k���,(nɽ�*<e����@��<�'!}��d��w����H
E#LPA�Y��gɽ�*<e��篐^������$�����~߿䳱`�t,\�����eɽ�*<e��C����.D.7�㸱�>c����]se���@=���r�c[�`t��NSad��ɽ�*<e��
���a޲�5����,ݞv�S��V
��u�3ba�d�ɽ�*<eP�7ٝGy�ɽ�*<ec�0�I7�ɽ�*<e�p�{��J�����cΔ_�`V�f�Bɽ�*<e����@��<�'!}��d��w����H
E#LPA�Y��gɽ�*<e��u<@B�*G���}�I#�L��~0H��r�dZɽ�*<ev���en�]�7�vE{��l��^5)��ɽ�*<eɽ�*<e�������1<�}���r�O�. ���ɽ�*<e��
���a޲�5����,ݞv�S��V
��u���*_ɽ�*<eP�7ٝGy�����p��S�\�(�|�C:���֌n]�0�����p��ɽ�*<e�̱Z︷�;�D`��G��Mc_�rɳ'ԙɽ�*<e�cǭ����d�S�F#)"cUm��Ȝ��X|�YA�Y��gɽ�*<e�q䆧K;y�0l�F�*���� 3���Z�
�A�Y��gɽ�*<e9�ݞR��=ɽ�*<e��ޢmo-e�;�Sx���]L�Eɽ�*<eƚ�������H��8�vE{��l��O�pٺe�ɽ�*<eɽ�*<e������;�3`-�}���r�O�. ���ɽ�*<e��
���a޲�5����,ݞv�S��V
��u�3�ӣR��ɽ�*<eP�7ٝGy�����p��S�\�(�|��4]���֌n]�0�����p��ɽ�*<e�̱Z︷�;�D`��G��Mc_�rɳ'ԙɽ�*<e�cǭ�����֘ڝ���x��F!Ȝ��X|�YB�<�k�qɽ�*<e:j���+�,�MG2˶��V1\�����s�>���K.ۗf��A�Y��gɽ�*<e�q䆧K;Jp�qKN�>k���,(nɽ�*<eɽ�*<e-H�x�kt�[~$�S��b�^ߣp�:�q>{=`b�D��t�[~$�S��b�^��ݵ�I�,O�`V�f�Bɽ�*<eɽ�*<e�p\�Ì����z�'Ɂ�}�����[3��f.�5i]΀ST����p��ɽ�*<eɽ�*<e�̱Z︷���n��U�0H��r�dZɽ�*<eɽ�*<ef�{��t�ɽ�*<eɽ�*<e�_F��x�������,�t�[~$����_��,��%����?Z�
��MMh84\Z��&���&S!i��g
x���]L�Eɽ�*<eɽ�*<e�يHc~���OX�gk�Δ�hYL�a⎣�S6��m���ɽ�*<eɽ�*<eƚ�������H��8�M�3pI^C�����p��ɽ�*<e'$��R��e�����kV�ɽ�*<eɽ�*<e}�tؤ�l�k���,(nɽ�*<eɽ�*<eܟ�	��ץ#�Xb�t�ɽ�*<eɽ�*<e��ɖ�Jb�ߞ3��㕵��\U+�;UI�&���.�Q�alZj2�IO����Z��\�ɽ�*<eɽ�*<eƚ�������H��8�ɽ�*<e{E�6��h#A�Y��gɽ�*<eɽ�*<e3%n�������U*��� a���!T��{%"��ɽ�*<eɽ�*<e������I�X��*�Å5�W����o�Ϗ��s��'�a?ɽ�*<e�P8񒽮ɽ�*<eɽ�*<e=���6���H� ȩ�꿲�~�~G9�!�Ҷa�c2U��<6|��V��@��5�ɽ�*<eɽ�*<e.�W�f�����ꖞ�Ж�x�3������t�7�P:�͎������(ɽ�*<eɽ�*<eO@�����w��d���cBGnň>�P���;�IzF}(hX�K��B=�Vz���.��Dd2vN���|�����p��ɽ�*<eɽ�*<e0�J���QWk�HZ�s��l�s��6�fz���Yr5ɽ�*<eɽ�*<e�6����iP��[P��x��F!���8�!�|ɽ�*<eɽ�*<e����,�4ɽ�*<eu:׈S�y|��5�L/%ɽ�*<e9�ݞR��=ɽ�*<ev=�H�U����ӯ�oM�\�l����������ɽ�*<eɽ�*<e��q�Ӭ�P�4�ׇ/�aU���ɽ�*<eɽ�*<e����@��l]AE��q�|�i41�����p��ɽ�*<eɽ�*<e��p^�S��	S&�4[�7������
:��{gɽ�*<eɽ�*<eɽ�*<eS�&��"x�R$��"�
�S�v>���GA9�n�@ɽ�*<eɽ�*<eɽ�*<e��E�5���s�!.�o���E�5���=��������
:��{gɽ�*<eɽ�*<eɽ�*<e�tR�\�5����<���^_��c�wF��b�Α��|�<78����Yr5ɽ�*<eɽ�*<ex��*��~�������ɽ�*<eɽ�*<e����@��<�'!}��#��T!uQ��NSad��ɽ�*<eɽ�*<eɽ�*<emk��畬��G��Mc_�rɳ'ԙɽ�*<eɽ�*<eɽ�*<e�9��w�[�����u�3���р�?���1�WNɽ�*<eɽ�*<e��8t������p��ɽ�*<eɽ�*<e�+�r��y�ɽ�*<eɽ�*<eO�
������$��5�yϦM�|.�`V�f�Bɽ�*<eɽ�*<eɽ�*<e��;��t��9.�0H��r�dZɽ�*<eɽ�*<e��8t������p��ɽ�*<eɽ�*<e���B6�]>����ueJ�1�	slEM�1�7"��ɽ�*<eɽ�*<eɽ�*<eL�Zo*̍��.��Z��X��7A��D	�)��)2���ɽ�*<eɽ�*<e���F5�K����'��S�K�n���oھi��͗
ɽ�*<eɽ�*<e2$6� 7�hx���]L�Eɽ�*<eɽ�*<eɽ�*<e3��h���!��ҳ�}���r�O�. ���ɽ�*<eɽ�*<eɽ�*<e���8o����^
�G��Mc_�rɳ'ԙɽ�*<eɽ�*<eu:׈S�y|��5�L/%ɽ�*<eɽ�*<et�ɳ)�Rx���]L�Eɽ�*<eɽ�*<eɽ�*<e3��h���!������1}���r�O�. ���ɽ�*<eɽ�*<eɽ�*<e���8o���31�y���G��Mc_�rɳ'ԙɽ�*<eɽ�*<eu:׈S�y|��5�L/%ɽ�*<eɽ�*<e�ag���x���]L�Eɽ�*<eɽ�*<eɽ�*<e3��h���!���r��qA}�U�V�O�. ���ɽ�*<eɽ�*<eɽ�*<e���8o�����+2j�G��Mc_�rɳ'ԙɽ�*<eɽ�*<eu:׈S�y|��5�L/%ɽ�*<eɽ�*<e|m�U!x���]L�Eɽ�*<eɽ�*<eɽ�*<e3��h���!g'�F5Y�}�U�V�O�. ���ɽ�*<eɽ�*<eɽ�*<e���8o��j3'Ƙl�,�G��Mc_�rɳ'ԙɽ�*<eɽ�*<eu:׈S�y|��5�L/%ɽ�*<eɽ�*<e'V>g�h�gƧ)����ɽ�*<e1��0ɽ�*<e����LT�D����x���]L�Eɽ�*<eɽ�*<eƚ�������H��8�M�3pI^C�����p��ɽ�*<eɽ�*<e����Xi��I#�L��~0H��r�dZɽ�*<eɽ�*<eO�
����8��i%�Uiy���mDx���]L�Eɽ�*<eɽ�*<eɽ�*<e_��B85���@z�Jɽ�*<eɽ�*<eɽ�*<e3%n�����%� ˙�ф�ӯ�oM�K���B6�ɽ�*<eɽ�*<e�&�|�D���}�ii��H
E#LPA�Y��gɽ�*<eɽ�*<e֪��"�+��bhF_����չ�<ɽ�*<eɽ�*<eɽ�*<e<�ʏG�ʓ�8�����G�Xz�(m{��v].����p��ɽ�*<eɽ�*<e�VJUT���[�a���`�?�B/�u�$H�-�d��\��Y0����Fb!�ɽ�*<eɽ�*<eɽ�*<e�cǭ���Ę(��I<�rPV��3�9�-���k[�*��m>6D��f��ɽ�*<eɽ�*<eɽ�*<e1��0ɽ�*<eɽ�*<e����@��js���JIa���P6x���]L�Eɽ�*<eɽ�*<eɽ�*<ewRۣB���n[�f�KvE{��l��^5)��ɽ�*<eɽ�*<eɽ�*<e�p\�Ì����z�'ɕ�R'�ސp"��˳c�ɽ�*<eɽ�*<eɽ�*<e,4���?w������7�5�.7���I{e�� �0��N��������JE���Dɽ�*<eɽ�*<eɽ�*<e�VJUT�����ޢ�CϮR�"d,!8�}�F@��ݤ�/���?�j�wyH'%Z��_.Fzɽ�*<eɽ�*<eɽ�*<eC!m�C���_ID�����Wre�	�&Ke�����E�����T̴U�ɽ�*<eɽ�*<eɽ�*<eO@�����w��d���cBGnň>�P���;�IzF}(hX�K��B=�Vz���.��Dd2vN���|�����p��ɽ�*<eɽ�*<eɽ�*<e5���.���'d�����I#�L��~0H��r�dZɽ�*<eɽ�*<eɽ�*<e�Y��#��Ֆ����E�ɽ�*<e�E��-ɽ�*<eɽ�*<eɽ�*<e�+�r��y�ɽ�*<eɽ�*<e��8t������p��'$��R��e�����kV�ɽ�*<e�jЛ4�1�b�R��x���]L�Eɽ�*<eɽ�*<eɽ�*<eZ��ފ�U�q<r�o�s���O����g�#w�����f�B��6�� Ɯ��g�#w��ٲAG������p��ɽ�*<eɽ�*<eO�
�������_2�'S��~�����)z��,sݻ���f�L5��	�.��,sݻ���f�&����ɽ�*<eɽ�*<eɽ�*<eZ��ފ�U�q<r�o�sU_��h�����g�#w�����f�B��6�� Ɯ��g�#w[��72�r����p��ɽ�*<eɽ�*<eO�
�������_2�'S��~��� �Lf!6Y,sݻ���f�L5��	�.���c5��I-�ɽ�*<eɽ�*<eɽ�*<e��ky�-��ɽ�*<es��l�s���
:��{gɽ�*<eɽ�*<eɽ�*<e\`/e�f�af�w��G��Mc__xZ��C�ɽ�*<eɽ�*<eɽ�*<e3M�ږ�ɽ�*<e��@�ї=D��}	��$?���1�WNɽ�*<e�+�r��y�ɽ�*<e�?���to�� a���!֌n]�0�����p��ɽ�*<eɽ�*<eC�=�%1�pі�_0g�ƛ����p��ɽ�*<eɽ�*<e4�0f2���W��#T������3�ɽ�*<eɽ�*<euQ }\�T�_.*=q�u�8tu�A=�t���y�Pɽ�*<eɽ�*<eɽ�*<e]�2T�A-��O�,�=/�[ٱ��@z�Jɽ�*<eɽ�*<eɽ�*<e�N�]�Kix�(͋Z�Ġ�mM�3pI^C�����p��ɽ�*<eɽ�*<e�ʚU$`�bF�1��;D
'��`�`3i��)�NSad��ɽ�*<eɽ�*<euQ }\���P�]��/q�u�8tu�A=�t���y�Pɽ�*<eɽ�*<eɽ�*<e9P�Ɣ���-��O�,�=/�[ٱ���-�8wɽ�*<eɽ�*<eɽ�*<eI�����8Kix�(͋Z�Ġ�m.2P:���[����p��ɽ�*<eɽ�*<e�ʚU$`MVR̤%);D
'��`�`3i��)C
�V[�ɽ�*<eɽ�*<euQ }\�x�}�@ķq�u�8t0φ8�	�tr*Nx �ɽ�*<eɽ�*<eɽ�*<eAx����'-��O�,�=/�[ٱ��1�,Wɽ�*<eɽ�*<eɽ�*<eW�VegW�Hu���~}Z�Ġ�m��s�P3�����p��ɽ�*<eɽ�*<e�����9�����p��ɽ�*<eɽ�*<eTϱ'���W��T�M�V�kCI�Ѣ��Y�8ɽ�*<eɽ�*<evS+ё@�Gܟ�ê.ɽ�*<e��B����ɽ�*<eɽ�*<e�VJUT���/�3�S�u��%e�܉��~Х���'�T ƶ�_��;ɽ�*<eɽ�*<e�VJUT������I�6lD������
�˦�2�RR(@��Ӯ�)��/�s�{ʪ�ET�,�:�ɽ�*<eɽ�*<e����n��r]���e�},�+���^?쮯���M�L>�;>c�)��kq��q�ow(������p��ɽ�*<eɽ�*<e:|Z�	����l�\�_E��Rۇ�d-�
��9qA�����xx���y�\7^��'^ɽ�*<eɽ�*<e,4���?w����p��ɽ�*<eɽ�*<e���4zm�
�K����Y�-B��, ��Ã����5�%j=ƚ�9����oS;������p��ɽ�*<eɽ�*<eȫ�$m4���Ɛ�����+e7�"��j3��aO������|G)�~�O��E������ɽ�*<eɽ�*<e�VJUT��ȭzE�'��v����Nހ��w���V`��1��zB7q@s�b2�M/��J��Yr5ɽ�*<eɽ�*<e���M����z�IYLy^�45R��K��/�žCɽ�*<eɽ�*<e��uf�O����OÞ���"'���A�Y��gɽ�*<eɽ�*<e.\��O����΄�ɽ�*<eɽ�*<eɽ�*<e��<��ݭ�`V�f�Bɽ�*<eɽ�*<eɽ�*<ee��Shq�M�L>�;>c�uۡ'��������ɽ�*<eɽ�*<eɽ�*<e����6��&��r�m�,[�+A�Y��gɽ�*<eɽ�*<eɽ�*<e7tO�M�Ͻ���8�!�|ɽ�*<eɽ�*<e'$��R��e�����kV�ɽ�*<eɽ�*<ef�{��t�ɽ�*<e��8t������p����-�e�/XM�Th ٞDw��s��JПE�[5ɽ�*<eɽ�*<e�i{ޝ��i#-Դ���Sk�k�9׎Oh���y��V�)iɽ�*<eɽ�*<e��}Gδ�-/���?��t<ŕV�(�x���]L�Eɽ�*<eɽ�*<eɽ�*<e����6��6�9b������ßɽ�*<eɽ�*<e��8t������p��'$��R��e�Ӈ�ɽ�*<e����p�����A!q���"'���֌n]�0�����p��ɽ�*<eɽ�*<e0�J�����4_�ڬt���y�Pɽ�*<eɽ�*<e.�W�f����T96M�3pI^C�����p��ɽ�*<eɽ�*<e����Do���װ�|�Bޛfe�^C�ɽ�*<eɽ�*<eɽ�*<e����tWn�]�7�M�3pI^C�����p��ɽ�*<eɽ�*<e.�W�f����T96�H
E#LPA�Y��gɽ�*<eɽ�*<e����,�4ɽ�*<eɽ�*<e���F5�K����'��S�K�n���oھi��͗
ɽ�*<eɽ�*<e�oc;�Eǎkn�f��H�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�#b;��3�P�^�#X7�I-��)�B�b� ��]�J��[�˒f�ɽ�*<eɽ�*<eɽ�*<e�Y��#���z�$�mj&�K>Z����-�8wɽ�*<eɽ�*<eɽ�*<ef�{��t�ɽ�*<eɽ�*<eɽ�*<e����^��	x���]L�Eɽ�*<eɽ�*<eɽ�*<e.�W�f��
�u��[��X����%Tϱ'���W��T�M�V��xX�-����p��ɽ�*<eɽ�*<eɽ�*<e�`��l�U �y1�P���R�.�����K��ǖ����p��ɽ�*<eɽ�*<eɽ�*<ed�p�c�-���x5���)�x)B[|,s�)5�RX�����p��ɽ�*<eɽ�*<e��8t������p��ɽ�*<eɽ�*<ea�E��x�.�`V�f�Bɽ�*<eɽ�*<eɽ�*<eO@����
/ ��Z��Z<�����,��w`&�j��~��Kn���8��#0A�Y��gɽ�*<eɽ�*<eɽ�*<e-H�x�k}^�R��R\wd�ԷD��K��ǖ����p��ɽ�*<eɽ�*<eɽ�*<ed�p�c�-���x5���)�x)B[|,D�1�	�����p��ɽ�*<eɽ�*<e��8t������p��ɽ�*<eɽ�*<eAjC����w.O��&x���]L�Eɽ�*<eɽ�*<eɽ�*<e.�W�f��
�u��[��X����%Tϱ'���W��T�M�V^�QW��ɽ�*<eɽ�*<eɽ�*<e<�ʏG���NIL�|T�"�ףG��T�A�Y��gɽ�*<eɽ�*<eɽ�*<e��؁�1��NILȭA�Ȩ>/Sc�>tFC�A�Y��gɽ�*<eɽ�*<eu:׈S�y|��5�L/%ɽ�*<eɽ�*<e'V>g�h�gƧ)����ɽ�*<eɽ�*<e{!�p�T**%w���
���g���ɽ�*<eɽ�*<e�يHc~�����'� ħ4��D T��)Y��W�ɽ�*<eP�7ٝGy�ɽ�*<e�i��c��ϧ4��D TT�D����x���]L�Eɽ�*<eɽ�*<eɽ�*<e�#ci�6�ɽ� K���+��pb5]\��~t�b�,�n��ɽ�*<eɽ�*<eC!m�C���_ID���s��l�s���
:��{gɽ�*<eɽ�*<eɽ�*<e\`/e�^|��]`�<��j_*��0���&��=�5K����^��C1"��L;D
'��`�Ϥ�^�	R�!�X~�h?�D��[)ɽ�*<eɽ�*<eɽ�*<emUF0�|���\'���Z�Ȱ����Z��XO���y�G$���=笥hɽ�*<eɽ�*<eɽ�*<e�pݰ
�g/���CvIO�:��E[=x<ݲa�_7ξkZ�x��`�])��ɽ�*<eɽ�*<eɽ�*<e? ѳ�ҵ
�ڝ�1�V�p��S	�����(���Ջ|2 kp�m`���JU�I+�ɽ�*<eɽ�*<e�VJUT����6���t�����gk�puLJ��8�{|�405C2V�����p��ɽ�*<eɽ�*<e�)�w׽�ɽ�*<eɽ�*<eɽ�*<es�����S��d}���{�hf��
�-A@78�/lI�Bdʓ}������ɽ�*<eɽ�*<eɽ�*<e<�ʏG����=�5K�0��I���/�žCɽ�*<eɽ�*<eɽ�*<e�d�ٝaAR[K�n��}	��$?���1�WNɽ�*<eɽ�*<e'$��R��eL�"۠��G���2�SY^!\�y�DpW�[x���]L�Eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�	��� �0�m!�]C��00�z�s��"/GP�vr�${˳ɽ�*<eɽ�*<eɽ�*<eɽ�*<e^��
�h���KI�"@HM��_{������3ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����O�02``4BFB1T���z���r�H��_�x�����p��ɽ�*<eɽ�*<e��8t������p��'$��R��e�����kV�ɽ�*<e����]��������`V�f�Bɽ�*<eɽ�*<e�VJUT���\��Ҧ�������3
���"�7R�f�D���9���0��N��~ɽ�*<eɽ�*<e4�K`��VR�w��d��#��k�2y���mDx���]L�Eɽ�*<eɽ�*<eɽ�*<e�`��l�U �y1�P��1l�XiI�����p��ɽ�*<eɽ�*<eɽ�*<e�9��w�[�s��l�sȴ��D��ɽ�*<eɽ�*<eɽ�*<e�Y�tѥE��䅓�g ������ɽ�*<eɽ�*<eɽ�*<e3%n����׿ȍ�rӭ�����m�ɽ�*<eɽ�*<eɽ�*<eP�7ٝGy�ɽ�*<eɽ�*<eɽ�*<e�r�_`�m��&�ӂ[uM�3pI^C�����p��ɽ�*<eɽ�*<e�+�r��y�ɽ�*<ef�{��t�ɽ�*<e'V>g�h�gƧ)����O�
��������H�GO4��F�̸B���l�Z)^��_������ɽ�*<e3M�ږ���le+�Ѝ�Ě��+����p��:j���+�݋��{��}���r�O�. ���ɽ�*<ewRۣB����G�O1�
��?�%�f�D���9��p���b�!�u:׈S�y|��5�L/%��"@�>���<��ݭ�`�*6Z�qD�F���Ҏ^0r��9��XM?s5n=E��Rx�5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��<�|j_����QC+��	�Uj�ǅF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��<�2��M]��()�8��q;8>�"��&A�}7g��q���9���,B�:��c �wRo�?��7���]� ��8���VP��͵@���o�?��7�1�h��HS��l�<ܺS^�J�Y�|���#2Ph�i!Mi���\$��N�<oJ;���}�^Cg5����q����c�ӳk��H��zw����C��&���Q�)y�
��2ˀFɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wF��M�C$#����p��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�0r�"��%����ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e:j���+�Y�\%�,� ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�Ɍ���%ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eC+��"=�t����m��cɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e"7�!ne*5�K\��t�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�s��"�w�[g�Ʊ�]ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eA�Jς��=����p��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<ecS�<�Uw�o��X ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e1Rk����`����p��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e`�!ܒ��]�������%�bR�xi53ة��Z����qp��Q�k��/�B��?;�{�ۥ�a\�X�}%�<�	�B�a�h�:׸d�9�+��_�i�q�k�אO@�������w�i�E�9����CI���i|���o��V6�B�a�h�"7�X�G�EA�:�W�.�^<�
:�:j���+��~�;5��\�I;���Ԋi4"�J�'{�0�79u��� ��#*ɽ�*<eM�T�9F�9�ψ���ɽ�*<e�U����7��̏W�Z������'$��R��e$1͉������Zɽ�*<e4��O�ջ�RKD�vQF�I6:\%X�(��j4�v�'��w4R�8�2Q�l-nL��^����w��;k��*Y�%^����͕��cW�7A݁���� Y8ڛ&���Ԫ�N��RN���Ȧk�v�����9��]�(������cW�``�vA�h1-��j��<ǅ O�����5ݱ�C��cvr��?u�X<z��'̕��cW��Vk_���;���#�����p�Y�|�h8׬6l:4Nb� 'o�^{(�0v��]�m�ʓ�-��&�8����΍��]27�G#���ɽ�*<e��c�ӳk��H��zw�|�>l���_"K��c����}G�����ٸ�ɽ�*<e�S�k�a�;à����uf��@�I�PӰ�oSC���ԕ��cW�f3���W���?��4�?�}h��=��(�
����H�6�YЮ����e�W�p\�Ì�Ep�+|�G���3O#Ey�뽬=T�%�ҥ#"������p���U� ��8U�6\FU4�cEs����XӅ��޷��þ���L�:�NQ���ɽ�*<e��.˼:Nn��txO�UԮ6�n�`��:��G}M���,�>�۫�i�u{9xɽ�*<e��L�Y��'o�^{(��T��5g�:��G}M���,�>�۫�i�u{9xɽ�*<e��L�Y��'o�^{(N��1��E���[��^I�|*�<A��mt�[(PD���_Q�'��yp�4�q`�����o�j\B�(�*=1`�ّ��0���E�M5׽�;N
RC h�4�ZC%�4��9k���j�Z���;N
RC h�4�ZC%�45ԛ��}�I��z�d� ���	O<�*1����9,εn��-��~	Q>���ě����qkb{٨� �
��OL��X�aҥ��b��*�~��Q�)y�
��2ˀFɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e(���٤r�!x"�#��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e���+�����cW�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�怦\wɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�f�P+tx;�l��xDɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e7��� h)��Rd�'�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�U�����GwE	�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�s��"�w�[g�Ʊ�]ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e:׸d�9�+y�2w��\�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e:� ���[=����p��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eX"��}ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e"4�R��׾(�f�2$�hb;��8�*���x1�A{E`��DF��t_(��Ow�:3X�]�n"��%Hd�g�q���W<:Kɽ�*<e��������0��9�5<�B�a�h�cS�<�U+3H<��׹�"�a �ǚ�ǧ�d9�ψ���ɽ�*<e���<���Vbd90a�N5�Dr��;8aȆ���7�m��p.�^<�
:�vS+ё@��k��\�I;���ɽ�*<e�&Z6[�ػN0B��wo�	h�[@۾}��i�U�&_�zN�����ɽ�*<e6)ܰnslRKD�vQFɽ�*<e6�T��~�՛ar��Z�.Zw��GV7�H2��XZI����Zɽ�*<eϜ�e�S(;��2��:7<�|D��o��-���B�%h�o�T��^@ҽΣ)8���M���b��P�2}2)҄gn��txO�U՘yӬ����8B`}��t�q��ɽ�*<eFLnV�4��M��Z�F�+��jd� M��<�ɽ�*<e�~sh��&+���l�`�ۭY��'�P��*�v�m+��)	�x��34;�[J�ҟ��:)��!Nl�s�NP��XP�զ(�iDk�(催w5���@Ԁ6U�-zkeYLu1Y��끆E�n)1Jf�kR������BN��fS���N?J����A���9׉�F��A����Ym�B�frb�����r�m�5ݱ�C��7������O_DK��:)Ɣէ套��p�Y�����Q��2O��v6�Ks��'����������1������YU��iS�+~FZјF����L�uQ�^hD�|'cl>o�Gx5��:tf����/_��p%wKSQ�
gE��;�����Ӕ�ȧ�b8V��p%wKSQ��F1�I�NtGw���,61�UZ�K�)���W��:
6f�B�dW��&��F���(�u�����9F|���C|�����N���Q�)y�
��2ˀFɽ�*<eɽ�*<eɽ�*<e!����Mβ�N� y�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eyR]�=�W�r!w�I%F�s[�'���06(�ɽ�*<eɽ�*<eɽ�*<e�7l&��F�+����v���z�� ���� p�������p��ɽ�*<eɽ�*<eɽ�*<e\���d!2v�)�y��¿4�T i���!�)ۂ%#Bɽ�*<eɽ�*<eɽ�*<e��_��l���]V&a;Bɽ�*<eɽ�*<eɽ�*<eɽ�*<e��Hѿc�ߔG�=��ɽ�*<eɽ�*<eɽ�*<e	�r�	�O%L�;?C��Oɽ�*<eɽ�*<eɽ�*<eɽ�*<eyR]�=�W�r!w�I%F�s[�'�5�vӸ=].ɽ�*<eɽ�*<eɽ�*<eɽ�*<eyR]�=�W�r!w�I%	�>zF, <�t-*����cW�ɽ�*<eɽ�*<eɽ�*<e�~�}����n2���/^��"������R���7�4�z�P�ɽ�*<eɽ�*<eɽ�*<eL��]�1#�A�E��W��NO��YWW��m!�~����R#l�J�Ǥz)J�.�;�Zi�I�wL��9����CI���i|��se]��.)����p�qA��=	oO�. ����eF9YH,ɽ�*<eyR]�=�W�r!w�I%	�>zF, <�t-*��0��9�5<�B�a�h��7l&��F�+����v���z�� ��#��k�2u�>��d�F��� ��#*ɽ�*<e@82�����9���z�4��Uv�p��v\H����.�^<�
:�kwO�&뿃_W��D����7R-��m�D��"�ەZ��K�N5�Dr��M[�'��
��p�N5�E��<)�a�8����O�. ���\�I;���ɽ�*<e�&Z6[�ػN0B��wo�	h�[]�����p�����RKD�vQF�I6:\%X�,+�)c�9���z�4��Uv�p���& �'��ar��Z�.ɽ�*<e\���d!2�\��'t:���:��DM�L>�;>c�初3�;Z������kwO�&뿃_W��D����7R-��R�q��Ң!�u�"J�4�2��R�ɽ�*<e���<���viI�$
���z!�l��;8aȆ�U����Z������'$��R��e$1͉������Zɽ�*<e4��O�ջ�RKD�vQF�I6:\%X1l��)B	�zN�����ɽ�*<e�QƖeK�RKD�vQFɽ�*<ew�ſ"h�Pa]��Ÿ��ch�c�y��UB}yh��꠰����Deϑ����>��>l��#�����T�/K��'�1����^ ��r��b��,E�E�b��i���sX!�_Өg%��5���]�H������ꡜ��|�J���ϲ\�I72�~sh��&+���l�`�ۭY��'�P��*�v�m+��)	^ ��r��b��,E�E�.=⨽9��8��d}��	�ё�uC�-��#�����������;v�88���í�2D)�<�e|��n��=�U6Ǉ0Y�U��ӻ^��|	g��i��@�r�y.���i�&�V�Zx���끆E�n�w�}{�D��"��`ޕ끆E�n]��ƚ����p��V�e���V�uCM꼤3_�}��Q����� D�x�J���#��xV��g���%�#�g�ަB qg�����6m<wm�;P(�Y�#lh�o�T��0��(/�� ��U�L>YJ�l�EOEM<C�)yR]�=��{i�x��U��l���;+���V��.>YJ�l�E&��E� ��t �)0�;\���'u���:��D͛���0�F��2Y�"e_W��D��w��d�K��H1�2Ϝ�g,��%�">YJ�l�E��ص'�D�t �)0�9���z�4��Uv�p���v��<����{���D"`꾶��~�;5��F��2Y�"e_W��D����7R-��R�q��Ң(H��u�6�C�-�m+*}��PjyR]�=�W�r!w�I%	�>zF, <�t-*�'A$橇�H-P�ġ|wug�Dp7�1X�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�d�D5Y��Z���5���&#�
�-%dC���sEU:�h�H�5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�^��'[�EE�}�^Cg5�<�]�=׺F��o������Ɯ�hm]�ɓ�tC"Ɔ�;��t�^	&2Bv�s��yl2���ɽ�*<e�G�x9��F�G��/�gj��� ��#*ɽ�*<e7��� hॗ�'#qݤ������a���D9$���$@���Ę�c5����_k`ɽ�*<e�C�.��MҼ��>i�5��M���>���6�����&B��E����Ѳ����{72L%hQQṏs�3(c]ǻ8_��&��!Q]���W<:K��{v���]�P�.�F"�#F��87U*���g���&B�����9��ɽ�*<ee&����h�V8��+ Zf�UgYavkF����{4�gvTM����n�Gl=�F��7 Z��6�*�ҵ{b��D�*��F���5�vӸ=].]�P�.�F�f�[>���ɽ�*<e*��F�����06(���� ��#*ɽ�*<e�r�_`�m��d�2I�n�ȳ��,h8���� ^��
�h_<9�I�E�ɽ�*<eةO�!�	/?�Ƹ��."x�֖�J��D��!��f>>_YRcy�q<r�o�s�<I��FM2��e��jɽ�*<e+�Ax �c��װ�|�B�d�'�_���4�t�ȧ��`�ȓ"`Õ�s�塰s�'�B|��;��KKɴ�3��l�?/��<�����K���*��q%'cX�Kɽ�*<e0�2���H�ʷ��� �9"�w���b"8��ɽ�*<eoP�}>]$��o����Z8�P��ؾg��t{2ۀHɽ�*<e4��؏���U=�j���k��V����U�zЕ&��|JПE�[5��L��$)�Q���75�w����ņ ���@��ZS��3�����kV� �ypC�G�]0;�G�	�M��)��3�uѨ�<��!����;��pY$x���]L�E����@��r�����cδ�C:Z���/�žCɽ�*<e�8z�z@�~��Kn��4�[�GC����|��ɽ�*<e���&B���ym��Aٰ���˫�M�3pI^C�����p��ɽ�*<ee&����h�V8��+ Z�G��Mc__xZ��C�ɽ�*<e��!�2X��..+`����x��F!��@z�Jɽ�*<e\Jԙ�% �f��S�Hɽ�*<e�`F����A�Y��gɽ�*<e3%n����ɽ�*<e�!TL�MUt���y�Pɽ�*<e.�W�f�Y��e�!�vE{��l��^5)��ɽ�*<eɽ�*<e,+�
����s�@��>�ڜ�O�����NSad��ɽ�*<e�nN�\�Rh{O�v;s��l�s����|��ɽ�*<eC!m�C��܍�P����>Է4M�3pI^C�����p��ɽ�*<e��;��t�c�#����G��Mc__xZ��C�ɽ�*<e�H)��k� mQ��5��x��F!���-�8wɽ�*<e�q�И�mJ��E|�m;ɽ�*<eɽ�*<e5&��j�Vހӝ3\x���]L�Eɽ�*<e\Jԙ�% ����'����V8��+ Z{E�6��h#A�Y��gɽ�*<e��!�2X��˃�6��Rb��uCdZ��@z�Jɽ�*<e'$��R��e�����kV�ɽ�*<e�.U�[�x�ɽ�*<e�'�$I��q,�}�����p��ɽ�*<e��3�ꭚ���Tk���,(nɽ�*<eɽ�*<eɽ�*<e5&��j�Vހӝ3\x���]L�Eɽ�*<eɽ�*<eɽ�*<e]�P�.�F"�#F��8#��U��Z{E�6��h#A�Y��gɽ�*<eɽ�*<eɽ�*<eKy�1�,��K�am@��z.�1Q��@z�Jɽ�*<eɽ�*<eɽ�*<e\Jԙ�% �>|
ϒ���ɽ�*<e�G��Mc__xZ��C�ɽ�*<eɽ�*<eɽ�*<e����tWn�]�7�ɽ�*<eM�3pI^C�����p��ɽ�*<eɽ�*<eɽ�*<e��;��t�c�#���s��l�s��\!����ɽ�*<eɽ�*<eɽ�*<e�]�~�%Bh@P��ɽ�*<eڜ�O�����NSad��ɽ�*<eɽ�*<eɽ�*<e�8z�z@"�d�;�vE{��l��^5)��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�קto�o�ɽ�*<e�I#�L��~0H��r�dZɽ�*<eɽ�*<eɽ�*<e�+�r��y�ɽ�*<eɽ�*<eɽ�*<e,��w�6�%ˮ����)�tBC�j�%~��$nnD�a���C��"'�c��9U-��[���Bɽ�*<eɽ�*<eɽ�*<e���5$�bȊ�~'q���kUD3QƢ�ɽ�*<eɽ�*<eɽ�*<eC!m�C��#izE�Y��x��F!���-�8wɽ�*<eɽ�*<eɽ�*<e\Jԙ�% �>|
ϒ���vE{��l��^5)��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e3M�ږ�ɽ�*<eJw��:���Q�g
���A�Y��gɽ�*<eɽ�*<eu:׈S�y|��5�L/%ɽ�*<eP�7ٝGy�ɽ�*<eɽ�*<e�����0$7"f�gtkn�f��H�ɽ�*<eɽ�*<eaТk嫆��-B��, �����)�8ɽ�*<eɽ�*<eɽ�*<eC!m�C��#izE�Yɽ�*<e��x��F!��@z�Jɽ�*<eɽ�*<eɽ�*<e�p\�Ì��	� ]�Mɽ�*<evE{��l�T���G���,[�+A�Y��gɽ�*<eP�7ٝGy�ɽ�*<eɽ�*<e�^�Q#�z�,[�+֌n]�0�����p��ɽ�*<eɽ�*<eɽ�*<eff��a{?R[��%�w/ɽ�*<e{E�6��h#A�Y��gɽ�*<eɽ�*<eɽ�*<e��u<@B�*G���}ɽ�*<e����%t��悹��c޶'1��Uɽ�*<eɽ�*<eɽ�*<eɽ�*<e�f ��.��NL���ɽ�*<e��;��1�W/���?��W�=P��'kɽ�*<eɽ�*<eɽ�*<e���&B����7zN-ɽ�*<e��x��F!�W�2�[N���Q�]���e�gܓ�ɽ�*<eɽ�*<eɽ�*<e.�W�f��
�u��[Q�ҡ���s��l�s�*��F����a������eV3HU�ɽ�*<eɽ�*<eɽ�*<e֪��"�+F��Yf{ɽ�*<es��l�s�*��F���M�J�xN��H�qɽ�*<eɽ�*<eɽ�*<e�����3t�b�Α�蓔'd������x��F!���-�8wɽ�*<eɽ�*<eɽ�*<e\Jԙ�% �>|
ϒ���ɽ�*<evE{��l��O�pٺe�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����p��ɽ�*<eɽ�*<eɽ�*<e���RJ�q��(m�'�,"��h�@
�_��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e a�\��$��P�6;7}$�T�1.*��F���U?�De�:���*���悹��c� �v�zO�9��Z(��`V�f�Bɽ�*<eɽ�*<eɽ�*<eɽ�*<e@9_@�R4�P2��V5�vE{��l��^5)��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e
1���P2��V5�ɽ�*<eM�3pI^C�����p��ɽ�*<eɽ�*<eɽ�*<e]�P�.�F"�#F��8#��U��Z�H
E#LPA�Y��gɽ�*<eɽ�*<eɽ�*<e���&B���V��P �޸����of�����Ro�C
�V[�ɽ�*<eɽ�*<eɽ�*<e�p\�Ì����z�'��m�A���gA�Y��gɽ�*<eɽ�*<eɽ�*<er�֏��9�y'Uq<B��B�Z�Y����H��0���<�I2%��P�6;7}4k�Amsxb��+OVJПE�[5ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��u<@B�*G���}��x��F!��@z�Jɽ�*<eɽ�*<eɽ�*<eɽ�*<e��S��fz.G5�td'���9���\�O�pٺe�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e^��
�h&ꬶ�Rɽ�*<eJw��:�������ßɽ�*<eɽ�*<eɽ�*<e��8t�֨��S��D{�S���-�V�����W���/�žCɽ�*<eɽ�*<eɽ�*<eC!m�C��܍�P����>Է4�G��Mc__xZ��C�ɽ�*<eɽ�*<eɽ�*<e\Jԙ�% ����'����V8��+ Z�I#�L��~0H��r�dZɽ�*<eɽ�*<eɽ�*<eɽ�*<e
����d�
�˦�2�RR(@��A�Y��gɽ�*<eɽ�*<eɽ�*<er�֏��9�y'Uq<B��B�Z�Y���������<�I2%��P�6;7}4k�Amsxb��+OVJПE�[5ɽ�*<eɽ�*<eɽ�*<eɽ�*<e���:��޿��> fK��x��F!��@z�Jɽ�*<eɽ�*<eɽ�*<eɽ�*<e��2� �p���<���^�S=������O�pٺe�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e^��
�h&ꬶ�Rɽ�*<eJw��:�������ßɽ�*<eɽ�*<eɽ�*<e��8t��}�tؤ�l�k���,(nɽ�*<eɽ�*<eɽ�*<eɽ�*<e3M�ږ�ɽ�*<ea�~��P���yAI>���xGʃ�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e1��0ɽ�*<eɽ�*<eɽ�*<eG��.s�xɽ�*<e'$��R��e�����kV�ɽ�*<e����[�oqM��		��q�w]x���]L�Eɽ�*<eɽ�*<eɽ�*<e�#�����j�<�U�q�G��Mc_�rɳ'ԙɽ�*<eɽ�*<eɽ�*<e�קto�o�ɽ�*<e�����Ro��NSad��ɽ�*<eɽ�*<e�J4�2�|ɽ�*<eɽ�*<eɽ�*<e��}Gδ�-Awo��o��� ,��I����p��ɽ�*<eɽ�*<eɽ�*<e�g?k�Vtև̸B���%{�����_xZ��C�ɽ�*<eɽ�*<eɽ�*<e��Y��1Ϫ�K��"������p��ɽ�*<eɽ�*<eɽ�*<e!�j�˪�Un�]�7��?�Y
X�H��@�Xcݪܱ��Kz���q��k���,(nɽ�*<eɽ�*<eɽ�*<eɽ�*<e
1���P2��V5��I#�L��~t���y�Pɽ�*<eɽ�*<eɽ�*<eɽ�*<e]�P�.�F�"vЅ\�6�Q� g���
:��{gɽ�*<eɽ�*<eɽ�*<eɽ�*<e��uf�OϠ���/J�F��x��F!$������#Y�a@��ɽ�*<eɽ�*<eɽ�*<ef�{��t�ɽ�*<eɽ�*<eɽ�*<e:j���+��������q<r�o�s�����3�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�?�tT���/�žCɽ�*<eɽ�*<eɽ�*<eɽ�*<e]�P�.�F��u�ǧ2�j�P�@k)���T�M�VKf�a��A�Y��gɽ�*<eɽ�*<eɽ�*<eɽ�*<e�+�r��y�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�ag���x���]L�Eɽ�*<eɽ�*<eɽ�*<eɽ�*<e\Jԙ�% �f��S�H��;��1�W�~��Kn�*����Ob��w�Eɽ�*<eɽ�*<eɽ�*<eɽ�*<e����,�4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e� mC��=�JПE�[5ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��l�G�䗎Ei�����)�B�b� �-�<�_>��w�Eɽ�*<eɽ�*<eɽ�*<eɽ�*<e����,�4ɽ�*<eɽ�*<eɽ�*<eɽ�*<eAjC���u�Mf��k���,(nɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��l�G��ɽ�*<e��;��1�W/���?���v�G�wɽ�*<eɽ�*<eɽ�*<eɽ�*<eu:׈S�y|��5�L/%ɽ�*<eɽ�*<eɽ�*<e'V>g�h�gƧ)����ɽ�*<eɽ�*<eɽ�*<e{!�p�T**%w���
: ���5�l�y��
R���-�8wɽ�*<eɽ�*<eɽ�*<e����@������H��@�Xcݪܱ��Kz"�?^̠���/�žCɽ�*<eɽ�*<eɽ�*<e�p\�Ì����z�'��m�A���gA�Y��gɽ�*<eɽ�*<eɽ�*<er�֏��9��W8 �+N�����p��ɽ�*<eɽ�*<eɽ�*<e�يHc~���3I�.�$�ÀϚ?���)��#���ɽ�*<eɽ�*<eɽ�*<e'$��R��e�����kV�ɽ�*<eɽ�*<e'$��R��e�����kV�ɽ�*<e��8t������p��ɽ�*<e�����9�����p��f�{��t�UoZ*M��A��mt�[�b=�D2�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�]^�h���ÿ�7:��wA��W���4|�(�K��1�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��8�:o��"����ݸ8؋ֵ|�����N���Q�)yT�K._*�?-	��1XLם�A�<�-ZH�m�q��~��Wɽ�*<e���r�<���cW�\�I;���ɽ�*<e`ύ���#0�xy��?-	��1XLם�A�<�ކ��v��Yic��ݤ�����a3m����@����xw����Ę�c5����_k`ɽ�*<e둰�~�N!G���R����~��W"}�� I���O��xx�yN�F�8I5��Oh`�wo�	h�[����@���:��e
��F�����Ę�c5����_k`ɽ�*<e�*�S� V8��+ Zf�UgYavkF������!ڱ��Ճ5�M����F��7 Z��B�a�h�ɽ�*<eAwo��o�V[<Y7�0Ϣ���N���6����=���!�2X���=��c��v]�P�.�F�f�[>���]��2I&����l�G�䗕��cW��Kn�:Ou
����.��S��fz.G5�td'P�TT�Iic��ݤ�����a3m\Jԙ�% �G������r7U*���gHv@�����Uj+����0XP�9�<�C�a�6l����W<:K=�?���-1o�Z����\�?�5��Oh`�"�^�R`ot���X��1�k����{72L%hQQ��p��u��d+�2��y�����&B�����9��ɽ�*<e����.�+���&B�����9���-�?�L�r	[Fu�YJzh RL/A��5��M����Ve���P���e,��X������Ę�c5����_k`ɽ�*<e��z���"� ���j�F��7 Z��B�a�h�ɽ�*<e/���?��@���j�TJ���l�VUQ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q��F&��
`�ĕ�#G�:����ti<8=�yQaX�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)X��DF��t�h:��G%�D�*k�l82�8km���~U*�D��|F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�&���y���Vﵞ����o����O
e��H**�D��|F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8����.��Zݪ+i�]����G\�wMx��ޒ(W�	�n+�U�nr�������w��U)�՛C[���I�ʐ����Ezv�LD=c@�LT��~��!i��6�f��Q8&��x�$m��JYw�8�r�rz����&��ׁ�����`���ժ3]���w��J��*�D��|F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�&���y���P`�ܬ>���}�yU�	�KC��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�S�P��w�G|���X�34��>æ��`��6Z�Ւn���#�n���7�)�"Y|4,(r�p�V	#�3)��,�MG2˶�G�آp3�3p�N������~8�,(r�p�V	=ܾ���N[�ӣ�pgN�ʆQ'�y��~qT�Tϱ'���W��T�M�V��4ud��E�p��u��dwRۣB����|}J®N�ʆQ'�ɽ�*<e�H��|��_�9I��>�װ�|�B*���m�ʤ/5��k��>	�u���׳�D�u�[0������с*��*c��:��nB�r�rz���r�mCj���*������ѝ��c���wɽ�*<e1���CS�o�x��lPX��g��(�t�Ke�%zQɽ�*<e����#^�	Qu�;r�/�?���4��7�C�!#% ɽ�*<e����#^�	��Fl�qX?���4��t�Ke�%zQɽ�*<e��oj�L������ă$�f�Q"Om�7�C�!#% ɽ�*<e��oj�L�����uл���f�Q"Om�t�Ke�%zQɽ�*<e��oj�L���Cx���4����D�-�7�C�!#% ɽ�*<e��oj�L���q��̿���D�-�t�Ke�%zQɽ�*<eq�1�%`�iýf84�~�sW�7��R�FJ�����p��r�j�	��/3���р�
[JJ�������"�v+����p����-�e�/X\E�g��^�b`�砅I�6�U��)����p����-�e�/X�Va@�ZM�S�#��p��~7������p����-�e�/X"�`�}~vt�S�d蕴}3��3�	-����p����-�e�/XM�Th ٝ�	&F�`IY9�}�����p����-�e�/X�yAI>����v�K��F��i��1�����p����-�e�/X�yAI>����	&F�.x��y�|8�0͵�Fb�l�VUQ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q��=�%�>}6�֮Be�%c�^Od��X�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8����T%�g'�(�[�v��0�5*�"p�x^�����I�s|ִ!��>]����/J�!#�崵����옋F�W���ʟ���X}��;���s��Awo��o�x����&��̱Z︷�&�G�Zr��|}J®�qY~�,"�9u��夣�P1޸��ϝ<��Uצt��y4��"���JПE�[5��}Gδ�-�HYd����ޛfe�^C�ɽ�*<ewRۣB���n[�f�K��x��F!��@z�Jɽ�*<e��S��fz.G5�td'6�Q� g��\!����ɽ�*<eKy�1�,��K�am@�"RDn�fZ=t���y�Pɽ�*<e�#�����j�<�U�q�G��Mc__xZ��C�ɽ�*<e��l�G��ɽ�*<eڜ�O�����NSad��vS+ё@�Gܟ�ê.ɽ�*<e{E�6��h#A�Y��g�����>�QWk�HZ�ɽ�*<eM�3pI^C�����p��֪��"�+��bhF_vE{��l���x+,ɽ�*<e0������|�/��=1��x��F!d���m��ɽ�*<e���7	��l#�˴��56s��l�s����|��ɽ�*<e�6����iP��[P�!TL�MUt���y�Pɽ�*<eu-�!�J�ɽ�*<e��/���_xZ��C�ɽ�*<e&tb�~ҦR�c�#��ѱ����Ro��NSad��m��p�	��*k�n(
���>Է4{E�6��h#A�Y��g��uf�OϠ���/J�Fɽ�*<e����չ�<ɽ�*<eR:�sg�
K�n���o��x��F!���|��ɽ�*<eg�Jo�sl:�w�Y#�G��x��F!���|��ɽ�*<eZ��#1�R�!�X~�h+�����_xZ��C�ɽ�*<e� ��H�&4�OI�:�U�Z&\dt���y�P�Y�tѥE��䅓�g ������L�r��NB��As\(����)-:E�����չ�<��Yr5��
������3��;Q���"�+��/�žCɽ�*<e�g?k�Vtև̸B���%{�����_xZ��C�ɽ�*<eKy�1�,��K�am@�"RDn�fZ=t���y�Pɽ�*<e��)�������-�s��l�s��\!����ɽ�*<e����,�4ɽ�*<e��q�Ӭ�P�4�ׇ�\!����ɽ�*<e�ל
ϙ� ����@��
�E��d J\�K�g�[��6c�/ߔ�6�� Ɯ��g�#wc�+i0����N��"ɽ�*<ewp���	2Y�[�A����[�Xw^��5]���	�.��,sݻ���f���D�-�C
�V[�'$��R��eo�
�0�C����L�8j���	��y��6�� Ɯ��g�#wc�+i0��T�S�ɽ�*<ewp���	2Y�[�A��O05�j�Σ�5]���	�.��,sݻ���fX��g��(�,���ɽ�*<e�:�>�֖�9���Iɽ�*<e����:�֌n]�0�����p��ɽ�*<e��!�2X��..+`����x��F!��@z�Jɽ�*<eɽ�*<e��q�Ӭ=�u��OY�I#�L��~0H��r�dZɽ�*<ef�{��t�ɽ�*<e�p�{��J��dI�b��`V�f�Bɽ�*<eɽ�*<e��q�Ӭ=�u��OY�I#�L��~0H��r�dZɽ�*<eɽ�*<e���g�#w�'�S 5l�ڜ�O�����NSad��ɽ�*<e��
���a޲�5����,ݞv�S�����	������o��	ɽ�*<eP�7ٝGy�����p��S�\�(�|�B�&~�֌n]�0�����p��ɽ�*<ewRۣB���n[�f�K��x��F!���-�8wɽ�*<eɽ�*<ed2/�n�)�x)B[|,e���r�Z��u�i��ɽ�*<eɽ�*<e�6�����*�O-�KxgE.L$�z]U�b����_�Z"t�r�P�Чɽ�*<eɽ�*<eN��d=c]��o|��f����z�'�2����f��#�I(�ɽ�*<e���Ɔ��"ɽ�*<es����B8�ݣa{sr}JПE�[5ɽ�*<eɽ�*<e�̱Z︷�;�D`��G��Mc_�rɳ'ԙɽ�*<e�VJUT��ȯ*qNe�u?!=�C4/�2��g�����ɽ�*<e:j���+�X�K��B=�����B��T�T��	�xd��Si ��t���y�Pɽ�*<eɽ�*<e:�.�</Y8���{�k�&5����J��Mf�ɽ�*<eu:׈S�y|��5�L/%ɽ�*<e����p��S�\�(�|���KP�k֌n]�0�����p��ɽ�*<e�̱Z︷�;�D`��G��Mc_�rɳ'ԙɽ�*<e����tWn�]�7���x��F!���-�8wɽ�*<em��p�	��*k�n(
���>Է4{E�6��h#A�Y��gɽ�*<e:��8싄FmP&�����+�D�?�N�P��Vɽ�*<eɽ�*<e:�.�</Y8���{�k�&5�������v^q�ɽ�*<eu:׈S�yg��VD�ɽ�*<e��oj�L��w=��}�ྮ/�žCɽ�*<e~4�R�T�����Ӱ���s��l�s���
:��{gɽ�*<eL�r��NB�����j�۱`	�02jtz@L�A��V�)iɽ�*<e��}Gδ�-�o�c
����d���oj�L��kSG3�qfɽ�*<e�
�9����ɽ�*<e�p�{��J�5n��-‛�`V�f�Bɽ�*<e����@��<�'!}��d��w����H
E#LPA�Y��gɽ�*<e:��8싄F�U�R��c�+�D�?�N�P��Vɽ�*<eɽ�*<e:�.�</Y8���{�k�&5����H��-���ɽ�*<eu:׈S�yg��VD�ɽ�*<e��oj�L���:/cg��վ�/�žCɽ�*<e~4�R�T�����Ӱ���s��l�s���
:��{gɽ�*<eL�r��NB4��0Fi�S�?����tz@L�A�~�b���$�����p��ɽ�*<e��E�5���b�1̟-Ito�V9��'��x��^����sɽ�*<e��}Gδ�-�o�cJПE�[5ɽ�*<eɽ�*<e��}Gδ�-�)*�Qy	�F���g�9�"�[e���{��)*�Qy	�F���1K���<2S鋅$z����p��ɽ�*<eɽ�*<e����6��`�T�����O����Dc�Jr�JX�-�a��ɽ�*<eɽ�*<e~4�R�T��ި�q1�v����-�8wɽ�*<eɽ�*<e��8t������p��ɽ�*<e'$��R��eo�
�0�C��)*�Qy�{ʻ���4�����E{H��W�t��=���+O����|�ey*�����`V�f�Bɽ�*<eɽ�*<e�p\�Ì��-�Rٟ"z���0EN�a�"�˂7�kɽ�*<eɽ�*<e����@��<�'!}��#��T!uQ��NSad��ɽ�*<eɽ�*<e�+�r��y�ɽ�*<eɽ�*<ewp���	JПE�[5ɽ�*<eɽ�*<e,4���?w��B#rhoɽ�*<eɽ�*<eӏ��,���#ځD����c�\�Hefˢ�졻�!����%�����a�>5~zJzɽ�*<eɽ�*<e�p\�Ì����z�'ɑ��\��S;���w�,ɽ�*<eɽ�*<eɽ�*<e{M�y0��bm�B����.�>Ƒ�C
�V[�ɽ�*<eɽ�*<e���6*�H$����[�!�?�e�e����A�Y��gɽ�*<eɽ�*<e[����Eh�P�,&f0H��r�dZɽ�*<eɽ�*<ef>>_YRcy�q<r�o�sAB&QEWŦA�Y��gɽ�*<eɽ�*<e��q�Ӭ�P�4�ׇ�\!����ɽ�*<eɽ�*<eP�7ٝGy�ɽ�*<eɽ�*<e1��0ɽ�*<e�
�9����ɽ�*<e�p�{��J�,�a��(�8��p��k���,(nɽ�*<eɽ�*<ewRۣB����G�O1�
��t.�y�aɽ�*<eɽ�*<e��
���a޲�5���ޛfe�^C�ɽ�*<eɽ�*<eɽ�*<e�6����BP��#�,��x��0H��r�dZɽ�*<eɽ�*<e�VJUT����� �р���S���c8��̢}z)�Vt�ɽ�*<eɽ�*<eɽ�*<e,+�
����xu�Tv�,+�
����l�+�%6�l0H��r�dZɽ�*<eɽ�*<e����@��&���k�K�am@��Yҁ�37��q<r�o�s���O�����p��ɽ�*<eɽ�*<e��&�������p��ɽ�*<eɽ�*<e�&�|�D���}�ii��E��o��ɽ�*<eɽ�*<eɽ�*<e0������z��ݪ�O�pٺe�ɽ�*<eɽ�*<eɽ�*<e�يHc~���'d�����ծ�	��V"��˳c�ɽ�*<eɽ�*<eɽ�*<e�+�r��y�ɽ�*<eɽ�*<e��8t������p��ɽ�*<eɽ�*<e+teM�i��˃�6��Rb鍴\�&�)��/�žCɽ�*<eɽ�*<ev���en�]�7�.2P:���[����p��ɽ�*<eɽ�*<e�+�r��y�ɽ�*<eɽ�*<e����n��r�ӭ����kK���Q���j3�H��>m����ɽ�*<eɽ�*<ek~�l�W���ձa�Jm,ڣ8�Ya�,
!��������a!� ����[Y�ɽ�*<eɽ�*<e@�^�~=,+�
����.D�G�+8aɽ�*<eɽ�*<eɽ�*<eMW��o77����p��ɽ�*<eɽ�*<e��݇%����h����u�Ȝ��X|�YA�Y��gɽ�*<eɽ�*<e�]�~���b\	y`�k��������Iy�ɽ�*<eɽ�*<e'$��R��e�����kV�ɽ�*<eɽ�*<e� mC��=�JПE�[5ɽ�*<eɽ�*<eɽ�*<eo�wa��~�3�v,(��?��jZ�2�8�d�	��ɽ�*<eɽ�*<eɽ�*<eh��J6��Ɛm f^�8�I#�L��~A�Y��gɽ�*<eɽ�*<eP�7ٝGy�ɽ�*<eɽ�*<eɽ�*<e����Ca��/�žCɽ�*<eɽ�*<e"7�!ne*5^|��]`�c@s|x��tz@L�A��V�)iɽ�*<eɽ�*<eɽ�*<e���g�#w���
{���f&�Rk��ɽ�*<eɽ�*<eɽ�*<e�+�r��y�ɽ�*<eɽ�*<e�����kn�f��H�ɽ�*<eɽ�*<eɽ�*<e0��������Α�8?&�g�{����a�Iw�����p��ɽ�*<eɽ�*<e֪��"�+�2�M4p*��qE�26����D��aɽ�*<eɽ�*<eu:׈S�y|��5�L/%ɽ�*<eɽ�*<e'V>g�h�gƧ)����ɽ�*<e9�ݞR��=ɽ�*<e��n
�/�Dw��s��JПE�[5ɽ�*<eɽ�*<e�&�|�D���}�ii��E��o��ɽ�*<eɽ�*<e"7�!ne*5f�af�w������Ro�C
�V[�ɽ�*<eɽ�*<e���ð1�j��rq��&v
������/�žCɽ�*<eɽ�*<e�����>��4_�ڬt���y�Pɽ�*<eɽ�*<eɽ�*<e
����d�q�1�%`��4�cn-����p��ɽ�*<eɽ�*<ewRۣB����G�O1�
����Iy�ɽ�*<eɽ�*<eɽ�*<e���g�#w�� �w0	�NSad��ɽ�*<eɽ�*<e��
���@KY�~��pE��q�he��k���,(nɽ�*<eɽ�*<eɽ�*<e.F��f�=PC[�`]�R_X�&,)l=t�&{.��>��������p��ɽ�*<eɽ�*<ekwO�&뿃�h�����a<g�!<H~!��/"ˮSL�fr���]̅5<=ɽ�*<eɽ�*<eɽ�*<ef�{��t�ɽ�*<eɽ�*<eɽ�*<e�i88��C��װ�|�Bޛfe�^C�ɽ�*<eɽ�*<eɽ�*<e��uf�OϨ�H��j\E�g��^��j�ա{ɽ�*<eɽ�*<eɽ�*<e��!�2X�������d<�Yԁ���|���-�8wɽ�*<eɽ�*<eɽ�*<e]�P�.�F��u�ǧ2�C��lj,PP��
B���)0�7_�ɽ�*<eɽ�*<eɽ�*<e[����Eh�P�,&f0H��r�dZɽ�*<eɽ�*<eɽ�*<e2tB]$�H��@�Xc�
]��v�ɽ�*<eɽ�*<eɽ�*<e�&�|�D���}�ii�{E�6��h#A�Y��gɽ�*<eɽ�*<e��8t������p��ɽ�*<eɽ�*<e�+�r��y�ɽ�*<ef�{��t�ɽ�*<e�)�w׽�ɽ�*<e�����s�$H����G	m�pD{�������ɽ�*<eɽ�*<e[����Eh�P�,&f0H��r�dZɽ�*<eɽ�*<eO�
���� ��\bm�X��Z������ɽ�*<eɽ�*<e7�ϙ��&b����Ś@�P7a˾|����p��ɽ�*<eɽ�*<eY[v�_�MW��o77����p��ɽ�*<eɽ�*<eY[v�_��g��!^v�!�(I�,_��]�0H��r�dZɽ�*<eɽ�*<e�VJUT����
������~��\U�(�t��g5FSu{�=ӣ%�ϒ`�a��ɽ�*<eɽ�*<e�VJUT�����\�5��ɽ�*<eɽ�*<eɽ�*<e���d(�JПE�[5ɽ�*<eɽ�*<eɽ�*<e]�P�.�F��u�ǧ2�Cm�Ր�ιɽ�*<eɽ�*<eɽ�*<eP�7ٝGy�ɽ�*<eɽ�*<eɽ�*<e� mC��=�JПE�[5ɽ�*<eɽ�*<eɽ�*<e]�P�.�F��u�ǧ2�)�x)B[|,,-�ĸ�lɽ�*<eɽ�*<eɽ�*<e��8t������p��ɽ�*<eɽ�*<e+3A,>3tp�`V�f�Bɽ�*<eɽ�*<eɽ�*<e���&B���V��P ��Yԁ���|���-�8wɽ�*<eɽ�*<eɽ�*<e���&B��~��\U�(�A�Ȩ>/S�>Yy�ɽ�*<eɽ�*<eɽ�*<e��8t������p��ɽ�*<eɽ�*<ex�m���`��uF�Zr�x���]L�Eɽ�*<eɽ�*<e�VJUT����
������~��\U�(W$��;Gɽ�*<eɽ�*<eɽ�*<eNM{9q���g?k�Vtև̸B���%{�����_xZ��C�ɽ�*<eɽ�*<e,4���?w]�P�.�F�"vЅ\�6�Q� g��\!����ɽ�*<eɽ�*<eɽ�*<ef�{��t�ɽ�*<eɽ�*<eɽ�*<e'V>g�h�gƧ)����ɽ�*<eɽ�*<ef>>_YRcy�q<r�o�s�6䒉����q<r�o�s)��J�B��A�Y��gɽ�*<eɽ�*<eO�
�������_2�'S��~��g
��V������ɽ�*<eɽ�*<eɽ�*<e3M�ږ���$�=:�m1����}Eɽ�*<eɽ�*<eɽ�*<e[����Eh�P�,&ft���y�Pɽ�*<eɽ�*<eɽ�*<e1��0ɽ�*<eɽ�*<e'$��R��e��~�Nx��ɽ�*<e��uf�OϠ���/J�F�� w�8��1s5�A�Y��gɽ�*<eɽ�*<e����,�4ɽ�*<eP�7ٝGy�ɽ�*<e��ڈvV>���Qԁ1�	m�pD{�������ɽ�*<eɽ�*<e<[��C_s�b�Α��|�<78��	[Fu�YJzr"N���絁�����Д�٪,)9Џ�^�A�Y��gɽ�*<eɽ�*<e<[��C_s�b�Α��hu�v��`#	[Fu�YJzr"N���絁�����Д�٪,w��~QJ�A�Y��gɽ�*<eɽ�*<e<[��C_s�b�Α��}���T��	[Fu�YJzr"N���絁�����Д�٪,���.Қ��A�Y��gɽ�*<eɽ�*<e<[��C_s�b�Α��٧�1�	[Fu�YJzr"N���絁�����Д�٪,��(���mɽ�*<eɽ�*<e�CVE�OjN�W��#T�3�RR\���B?O榼W��#T��nb�~c�q<r�o�s��޶(:ɽ�*<eɽ�*<e(z�E%x �ɽ�*<e�I#�L��~A�Y��gɽ�*<eɽ�*<e3%n����ɽ�*<e�N�;�s3w���8Z�$��߁�Tɽ�*<ef�{��t�ɽ�*<e����[��"DП&���z���/�žCɽ�*<eɽ�*<eۓ]d�����~��Kn�Fj�g0��-�V���Аi�$��;ɽ�*<eɽ�*<e\Jԙ�% �f��S�Hɽ�*<e�w���xt!�Ж�x�3�A�Y��gɽ�*<eɽ�*<e��$�͛�ɽ�*<eQ��l(����Yr5ɽ�*<eɽ�*<e�����c5/���?��-���:�mc�� �@��g����Yr5ɽ�*<eɽ�*<e�Gx��y���6���́ZЍC0�v��U=�j�Q�����p�V'*⭦�[�轰�N�ɽ�*<eɽ�*<eɽ�*<e`s�����в/�M�	c�n�����s���W�%?�"��ra�%z(9YCQ��*����ɽ�*<eɽ�*<eg��xK�>5��
�殃3�:���&-��MsY|PD8���ԓ���iEz$b>W�����p��ɽ�*<eɽ�*<e���HGɽ�*<eɽ�*<e�/���g/�j�d�F�gc[�{�pj�~+yZ�H��=��>[�X��s�������ɽ�*<eɽ�*<e�#���;vf�c�����)*�Qy�o�\�Ҥ�E�,f`�V@�R����VG�g~#|��5�L/%ɽ�*<eɽ�*<e�Gx��y����}K�%)�X�<#��Rw�3�{Q�ۂ�0���z�IYLyh�t�E��ɽ�*<eɽ�*<eO�
�������O�U�!�9�y�E�JПE�[5ɽ�*<eɽ�*<eɽ�*<e����6���������)If�����tɽ�*<eɽ�*<e�i{ޝ��i�V�F\Z����p��ɽ�*<eɽ�*<e�q�И�mJ��E|�m;ɽ�*<eɽ�*<eɽ�*<e���ð1�j��rq��&v
������/�žCɽ�*<eɽ�*<eɽ�*<e3%n����׿ȍ�rӭ)�X�<#�?���1�WNɽ�*<eɽ�*<eɽ�*<eo0�ڝ*����g���ɽ�*<eɽ�*<eɽ�*<e1��0ɽ�*<eɽ�*<eP�7ٝGy�ɽ�*<eu:׈S�y|��5�L/%ɽ�*<e����Nހ�ky�Y��H�`V�f�Bɽ�*<eɽ�*<evS+ё@�ab��Z<�����,�w���xt!���$�O�
�w�Eɽ�*<eɽ�*<e���6*�H$��b��M&"_`���a�-�V���gڄ���ɽ�*<eɽ�*<e��
���ׂƯ78������h���`V�f�Bɽ�*<eɽ�*<eɽ�*<e�d�ٝa��@�ї=D�U=�j��D�B��ɽ�*<eɽ�*<e��8t������p��'$��R��e�����kV�ɽ�*<e
�˦�2�RR(@��֌n]�0�����p��ɽ�*<eɽ�*<e�#�����t,�a�¿�rɳ'ԙɽ�*<eɽ�*<e��!�2X�������d<�Yԁ���|�'l�X�.ɽ�*<eɽ�*<e���&B���V��P �޸����of
]��v�ɽ�*<eɽ�*<eɽ�*<e2Y�[�A��O05�j��ޛfe�^C�ɽ�*<eɽ�*<eɽ�*<e��2� �p���<���^%{������rɳ'ԙɽ�*<eɽ�*<eT��%z�����p��ɽ�*<eɽ�*<e����Do���װ�|�Bޛfe�^C�ɽ�*<eɽ�*<eɽ�*<e@9_@�R4<y��Ѹ@5�^5)��ɽ�*<eɽ�*<eɽ�*<e��S��fz.G5�td'6�Q� g���
:��{gɽ�*<eɽ�*<eu:׈S�y|��5�L/%ɽ�*<eɽ�*<e@�^�~=,+�
����.D�G�+8aɽ�*<eɽ�*<eɽ�*<e=����u�����p��ɽ�*<eɽ�*<e���&B����7zN-��x��F!Tϱ'���W��T�M�VKf�a��A�Y��gɽ�*<eɽ�*<eP�7ٝGy�ɽ�*<eɽ�*<eɽ�*<e����Ca��/�žCɽ�*<eɽ�*<eɽ�*<e��l�G��ɽ�*<e��w`&�j��~��Kn�*����Ob��w�Eɽ�*<eɽ�*<e��8t������p��ɽ�*<eɽ�*<e:<��f��k���,(nɽ�*<eɽ�*<eɽ�*<e���x���,49�iv (#X7�I-��)�B�b� �-�<�_>��w�Eɽ�*<eɽ�*<e��8t������p��ɽ�*<eɽ�*<eW�VegW��r�-�?������ɽ�*<eɽ�*<e\Jԙ�% �f��S�HvE{��lҵ~ԫ��G�&'hK��aɽ�*<eɽ�*<e'$��R��e�����kV�ɽ�*<eɽ�*<em{t�_�ͼ�(�nf�ɽ�*<eɽ�*<e�d�ٝa��@�ї=D����'������3ɽ�*<e����,�4ɽ�*<e4��؏������'�&���z���/�žCɽ�*<eɽ�*<e��)�����s%��r���
:��{gɽ�*<eɽ�*<e��
������3��;Q���"�+��/�žCɽ�*<eɽ�*<e��#2M)���x5���)�x)B[|,��D�����p��ɽ�*<eɽ�*<eR:�sg�
K�n���o�>��{f�CK�n���o��xt�%������p��ɽ�*<eɽ�*<e��!�2X���X"��|���@z�Jɽ�*<eɽ�*<eɽ�*<ejc)k�(X�,w/b�=��QGH�K�k|�����^#z�R�au���Mɽ�*<eɽ�*<eɽ�*<e�pݰ
�g/���CvIO�:��E[=x<ݲa�_7ξkZ�x��`�])��ɽ�*<eɽ�*<eɽ�*<e݃��V[�Ь�)x��_	�6���$�9Q.�G�/�.��{�7�?��|��5�L/%ɽ�*<eɽ�*<e����n��r�M_��[��,�X7A�@E��V�Zace��5��hi%��ɽ�*<eɽ�*<eɽ�*<e�ל
ϙ� ɽ�*<eɽ�*<e,4���?w�C�)ʹwW^#z�R�au�ƺf�L�����Ick]�x���ӇG����ɽ�*<eɽ�*<e��
���X�F:Ay���(#j��JПE�[5ɽ�*<eɽ�*<eɽ�*<e^��
�h���Q2�^�1����}Eɽ�*<eɽ�*<e�VJUT���R��^~���E�5���5��� *��k��M#���]Surw�Oc���y�G$����p��ɽ�*<eɽ�*<erL۪w�Ibk���g��H��#3���jЛ4�����L��hɽ�*<eɽ�*<eɽ�*<e��<��ݭZ��ފ�U�q<r�o�s���O�JПE�[5ɽ�*<eɽ�*<eɽ�*<e��}Gδ�-C-T ��>w���I�i����A������ɽ�*<eɽ�*<eɽ�*<e��^��t+���Er�y���:��`h�.i�t�ll�\&e��0��N��~ɽ�*<eɽ�*<eɽ�*<e���7	��l����7���eX����UU�im�aɮ��mF#[��A�ɽ�*<eɽ�*<eɽ�*<e����,�4ɽ�*<eɽ�*<eɽ�*<e^��
�h���Q2�^����oI�-6A�Y��gɽ�*<eɽ�*<e����n��rM���6�@���
2z?zo��E�5��ܶ���2v�-ɽ�*<eɽ�*<eɽ�*<e�q�И�mJ��E|�m;ɽ�*<eɽ�*<eɽ�*<e��uf�OϨ�H��j�yAI>���xGʃ�ɽ�*<eɽ�*<eɽ�*<ef�{��t�ɽ�*<eɽ�*<eɽ�*<e�ʵ�� Y��,�[m�}�ii�9��������5��1R	��B~d�x����B `8ɽ�*<eɽ�*<e�VJUT����b�vTP���m�Ƒ�ɽ�*<eɽ�*<eT��%z�����p��'$��R��e�����kV�u:׈S�y�R/�P�ɽ�*<e���5$�b��c�O��85"�#F��8U�v��<ϬJПE�[5ɽ�*<e^��
�h�&5���|��h���ɽ�*<e��#2M)��9/{��*ɽ�*<etz@L�A��V�)iɽ�*<e��q�Ӭ�P�4�ׇ��
:��{gɽ�*<e�+�r��y��X�OcB�+��p4�n��0��r�pB:�zMzՋh/Zk���kh�q}Rk!��^�(
P�����b�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�<Qs��'R?��9~�	��`,D��Y�0��s���M����飳������?ʌ�of�F�].���$��Jy�#@�����N�,9�{M���)_d<�cYb�'����4�È}����Hc�;�Y^�U=���8��u��(�H���-)�|�d!d�H�d�h�ݔ�x��{��õv�̟��������.s����g ��$�Lr�S��������N����!6���f����!Lؒ&�bL�.��. ����lB��,zyj���0_��A�\��B� �f����?���wIF�	D�$�=UQQ*rbH�iA�UAKTnО�>����x�})I)���()�6��9w2sO@�O�lK���K)��F��P���I1�3�䋇�æ��tg������a��4W%��g���$�-�����L}eW�+���{T��qɮ��B���(���%��|`ଽ��p�N_�qe�
��bS�����"�N�?�����LV7�q�BH�������(�k�T���cD�HM��נ#s��3��.5�)(�/��>4���3��h1��.�֊VG/"���@V��"W���à\j����f���ԝh<Kaչ�z�Mf%�l�J�����7N?����&8Y�`|X�+�2
���������h�>K	�K�7	�j����m%p7m�R���|"ÝW�qe�
��S$�����s�SŠ��z��Qd_No��t��C��[���d�bl�uxK|q�Y`h��1�D���_�2UE<�f��p'��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�/I�T���cψ5����4���m.o}��y���p%wKSQ��F1�I��}(��گ8�:o������4\���鳣���`��V�,�W]�ͻlU���(�����-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�)V ٥�Dk�͝�b�֏�V����5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^��DF��t��KJXx ��C��z��.d�)Qg��ϧ�p~rև�C�L��-<��eh�V��0�Bc��\�u�<T_����Zy=;��|�J���ɽ�*<e�6 �� |���DF��t���0UH�i7|2d>7E��O���"�*f��p~rև�
���F"xL��+�
"-w��-\�u�<T_2��G�= �B���R��bT�>Hw^���]��������mA����K��q�-�m�z_fN�d��t=X��Q�k��/޹���w쑣�gW�Yi}�_CQ>M,�Q�.#��W*͓M1�@ͫ�����e�ʝHw^���]�������淛}ذ�� �.�A�}�#��=:�mc�����F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)X��8ԟA��qO�싱�${��\yUL�4�v�Dm�b��Z��XO3΢B,�%,|,:�@vF�A�#u���^��?
�(�5��_��R���]��q5���E YPk�����xHL�ޫ
��U�61��Ţ/�ܻ�{X@��W�x���	�P���N��g�kq��;���S��TQ���=����[����o���5l�H����~�9�

?����HG�8���a*Ze���3;��ҩC3b\E��"Ϲ�t�:�e)(Q@S�6����W$cN7躜ȑզ�WH�&�ܠ��)�/������Һ��`h�X����Ft
��4`i
�8��W��/�ܻ�{e�T������������1���!�qHy��[���q�Q���\����� At�'� �dew�q�I�3O�_#g5�w�2����ey_6i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q��]��������7�e�;��X���2� �ߕ�"���t=X��Q�k��/�Nӹqs�<$�l=�F�=���qS-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�)V ٥�DkL�@���ڙ2�<;ۍ�	�:����8�����F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)XM,�Q�.#��e�x��W��b!�݊`�ͻ�8�g���=
�r�%�K!�R�Ժ�U@ͫN�)M,�Q�.#�R~�r����F�y���z�,U�n[��4N��� ��C��z��%�E �N���.�g{kX�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�T�N�:Y�?1�d�4D`�YZ͆ˎ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��o���ٽ�5����_k`ɽ�*<eɽ�*<e�l��m	5��Oh`�wo�	h�[ɽ�*<eɽ�*<e��^O�f5��Oh`�����\��.ȯY����Y��`#^��qQ0G]�Ҽ�w	�B�a�h�ɽ�*<eɽ�*<e�x[���K&���>��y~5����_k`ɽ�*<eɽ�*<e<�M��E�!�(I�=LU[$"��� ��#*ɽ�*<eɽ�*<eƚ�����˃�6��Rb=LU[$"��G�P�!����	*�sI���:Oژ�3�>������/�ĕ���KOM����(n�3y���]�Ҽ�w	$�.�prǿ8s6��Zv7��,�$��#B������6s�h$U+����.`s宍����w������G�P�!j9��y_ϰ���KK&���G�yB=�u�@3��6s�h$�d�_��wc���ġ}�3ě����6?���:�ɽ�*<eɽ�*<e~4�R�T��r{@ �P�G���W<:K� �h��ӟ�H�qҺ<[�������FaȫһAmic��ݤ�����a3mɽ�*<eɽ�*<e91��?��o8{��w��6?���:�ɽ�*<eɽ�*<e��S��fz.G5�td'P�TT�I���W<:Kɽ�*<eɽ�*<e���&B���V��P ��s��7Z�5��M��̦\;,N1f(��F�y���ң�:�C�Ť�ɡp�Z�Z8`���:��$uZ�i��9{y�2w��\�h�!��q��i��C�I���:O�g)â���ޫ�*�������*��dtKb����|ٲM��1���ۜ��G�~�L���㜗���d��̇�3͸8yw�T�+	4���Dg$ ې�b> |�!N5��Oh`�wo�	h�[ɽ�*<eɽ�*<eAwo��o��c�e[�J�VF�N4������w쑣�gW�Yi3Ȣ���o�ҳ�mxS�:�ug;
s郝��ɕyl2���ɽ�*<eɽ�*<e:j���+��Y�f�.��"�����.�^<�
:�ɽ�*<eɽ�*<e��\�����j�j�+��]���K-�c�g��*Kvɽ�*<e��b���i���!�)�0�s[+�"�72L%hQQ�տ�PK���)-:E����CW_s���1�k�eM�z{�����fם$�:Z������ɽ�*<e	H_0��J�����'���&��!Q]�eF9YH,����Zɽ�*<e�6�/��T�Xȡ�m��/���
0C���>MX�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�T�N�:Y�?H?cu���͝�b�֏�V����5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^x\��斳q4I�\6�0��<��f����J1.���d�Qd�����;xc&z�j��S�#�����d":r���4GHF�+��jd�ARË����ow����b�L:��X_��L�H��i]J�"䀊��� ]2&��4�H p~�rj�*���Nq�0a�L��+�
}�M���Qv��J��X��f������p��ɽ�*<eHc,�L) b����z�#d��!��f*��_�<v�z�u��Z ��Rji��p�ނ��:�.��zɽ�*<eɽ�*<e!��ɭK����é��U���#B����u�2��] yB=�u�@3~�=�F�GC��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S���������A�8�X�3VU=f�:>-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��m 	���`[�qW{���2I���)��Q��14%FD_�	�H"b��2W�T�m,�ZVG3���X�Mة>�w�~�d0Xl�5�����v����3#:%� 2]����j1� ^j�!ZVG3����B�X�Mة�*�����LA�Փ��H�iz�_d�Ar�3&�GE��7ۅ���z�%̗�Xl�5�������]4��<*�o�N�
�I���+W�L�q��� E�����&1�Rw�1w+>@�� Z(`���8�W�ޫ�*���,uX����s
�ڝ�1�V	�	n$�n�@�� Z(`���8�W�ޫ�*���,uX����s
�ڝ�1�V�\,��jΣ��g���ӅT���9�<Ѻ�w�u��V|��s�Ɂy����H��U�H���4�x3:Gv��S�P.�Y�S��:{�Z�'���I��zD��mJa�*��N���ú]'E���iO��А���
S�B�C�=�p?i@����Zm��02-�N�A��� Xl�5�����O��xx@^k-�Τ�'wL��͠�?�Vl��n��â����~wo����Q�wŋ���
�f=r���Ⲧ��b��.q$�A)�^U��얰�s��q��� E��mJ���M*� ���X�MةN��˅����w�TZVG3�����G���`���t�x�x�1��2��N�ʆQ'У얰�s��q��� E�	CI��X��q)
���"��m�
9r�)Q����v^����|��.E��7ۅ��e��O��&�!e��R���F��{�N�ʆQ'Щ�ѪM��u~�y‮��>j!aލ�\g��qX�Mة�A��G�|
[�:'�\�(�=�O%�o2����2I���¶���Xl�5���Q���c���W���gE���8�!�|��ӅT���9�<Ѻ�w�u��V|�oS�&�^�L�����]'E���i��D-	H_0����Iv4�4�z>�H4�'���2I�����h#Py�]�Ɵ�l�~�«V���34��1YϠ��.nx���qg+߄Fdd�r��H�;]�֙$D�ŭ�}�_�w��#ӡu�3l3I�}�2�aF�N�ʆQ'�ɽ�*<er��Ja����(�g�;vV��ؖ�8�u
����.A ɗt1$]�r��oR*lZAu
����.��G�H�BD�V���(d^��a�^���jJԔɽ�*<e̈�!��3�������z�8d�Gu
����..�W�f�X{�YyBҢ��s���N�ʆQ'�ɽ�*<e���cT�Bq�w��CX�Mة�p��u��d�.C��,����d��0���5���RKD�vQF"7�!ne*5.�z͵�$V���34��1YϠ�u
����.��G�H�B�U1��T+�A)�^U�ɽ�*<efE�4��^�)]%�CF�A)�^U�ɽ�*<eg��n6��RT��z6o��?�Vl��nɽ�*<eo0&%fw����F%�dC����yRKD�vQF\Jԙ�% ��/[-��!z:j�^�St�ar��Z�.ɽ�*<e��P'�8O�SH���͛ar��Z�.ɽ�*<eo�BUzZч-���ar��Z�.ɽ�*<e�*E��: � -�+�A)�^U�ɽ�*<e�(�ٮ@X{C����E��7ۅ��&ꬶ�RO�2�	��ǳ�y�|:j�^�St��{v������I�B�R�
!�ŮmaaU~Ξ�4N�ʆQ'�ɽ�*<e���>j!aލ�\g��q��Y�
D�I���jV���34�"��m�
9�5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^7�V<�N����X(-זauQ�s9���S��D�jCd�w,{� ��ps�g�nf3�g@����U1���]z/iq��{�9!��I��a|�k�e����H$k^��t���CE��d׽�-�~�}s$I����Q; ϋ5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^k2�G�CzӇG�����Z��
�Ť�ɡp��Z��uq:��GB���믏]Ep�����p���j�8]����ס����Ⲧ�2Xo�못oL��D�h��m�B����7��gt�K�am@�M�Fd�����r@�*�ɽ�*<e}��Pj�sɅ����!�(I��*�eM�[M�"vЅ\�����4��	s�o#q����tѹ�Ⲧ��b��.q$'$��R��efǢ�ڙ �.�Qq�*d��PtD���K>3���x��#e5�ɽ�*<e�(�[�v���~����(��MZ�/�y���!C�ɽ�*<e��^/a��헃P�� ��_�Iu��fz3:�(���V8��+ Z7L�XҪ��V8��+ ZyO$�,�cekwO�&뿃"^ym�4׼��'����V8��+ Z��t�H��,�K�am@�; ��?r��O�u��	F"B6�����p���+�r��y�����0b��*��-`�k2�G�CzӇG����%�hP��Fj>· ����	�N%� ���N�9Dݺ��ɽ�*<e����Ol!!��H/������K��8v�u>) ��`<�ɽ�*<e����@���e����>J͸8yw�T�����K��8v�u>) �]j�Q��ɽ�*<eɽ�*<e�(�[�v��^9�\ߏe�6VN�9� ����&��|l��I JF�7�\��F��q~�1"�ۻZ����K�`yO$�,�ceɽ�*<ekwO�&뿃"^ym�4�t�e&5�w�|l��I ������?BDiAx��E�^Ĩ�1��)�7h������_ԛ\�H
��x3:Gvɽ�*<eP�7ٝGy�ɽ�*<eɽ�*<e���g�q\i�>J����B�S�R#��(�nf�ɽ�*<ekwO�&뿃�`��$N��M�U�帶�<�+q�@J�F+�m9Kɽ�*<eɽ�*<e��^/a��헃P�� �9�t& �Τ�}��:+#�{�yPn;�ư�(��v��焄�D�#Gɽ�*<eɽ�*<e��^/a÷�&S)�
:@^k-�Τ��}S=:�����l�G���@RC��#L@=���\�H
��x3:Gvɽ�*<eP�7ٝGy�ɽ�*<eP�7ٝGy�ɽ�*<e �.�Qq�*d��PtD���K>3��Ĳ�<χ/�ɽ�*<ekwO�&뿃�`��$N��V����2��<۵!��,�[�>i �ɽ�*<e��}Gδ�->R}9�����k%J�?1l�XiI����� ����{��"�ɽ�*<eɽ�*<e��x�h�2��B������Vz�,@^k-�Τ��}S=:���#^��qQ0GB����3�����F���ɽ�*<eɽ�*<e}��Pjq��^U����_�Iu�� ⟒��d����%0)�7h������_ԛ\�H
��x3:Gvɽ�*<eP�7ٝGy�ɽ�*<eɽ�*<e���g�q\i�>J���d��� ��(�nf�ɽ�*<ekwO�&뿃�`��$N��M�U�帶�<�+q�@J�F+�m9Kɽ�*<eɽ�*<e��^/a��헃P�� �9�t& �Τ�}��:+#�{�yPn;�ư�Q�����<ɽ�*<eɽ�*<e}��Pjq��^U����_�Iu�� ⟒������"[���0��x�1��2��ɽ�*<e'$��R��e�����kV�'$��R��e�����kV�f�{��t�'$��R��e��䅓�g � ���N~+�{*9gƧ)����(��Î�HX�m��c\Nr��O�u�M�(�bJR���g���ɽ�*<e����Ol!!��H/������K��8v�u>) 9���
� �ɽ�*<e����@���e����>J͸8yw�T�����K��8v�u>) �l�JO�mɽ�*<eɽ�*<e�(�[�v��^9�\ߏe�6VN�9�#^��qQ0GM�����9�//[d���5��ӌfɽ�*<eɽ�*<e��^/a÷�&S)�
:wٵzfX����|ٲN��p޴o��o�s�,��2�0����Z�!�ɽ�*<e��8t������p��ɽ�*<e}�tؤ�lڠ8v�u>) g�3%�U877�P��ɽ�*<eɽ�*<e�Bk��٩1�o%��	o;�d�|�݁��!8����p��ɽ�*<e�j�8]����ס����9��@�Ixєf�,;��=VP����<hɽ�*<eɽ�*<e}��PjI�/��A�W�� 奫h(��2˲M@.F�rqD74�����ɽ�*<eu:׈S�y|��5�L/%u:׈S�y|��5�L/%�ŕI�(^�W8 �+N����� ��x���S۸����p��ɽ�*<e�����Q��/1lG%��,j˟W�ч-��ɽ�*<e��
������ ���7e���5��ri�`��i�>J���_��Bɽ�*<eɽ�*<e}��Pj���Mu���bZe-�q��+�ى�7�ϰ1�d��_��'D}��ɽ�*<eɽ�*<e�����Q����l��IŬ�!;,5�	/M7A���0��x�1��2��ɽ�*<e'$��R��e�����kV�ɽ�*<ewp���	��GB���X�0֊�Ն[�e����ɽ�*<eɽ�*<e}��PjN��p޴��B�)��c���ġ+CǺ�Q��ɽ�*<ekwO�&뿃����w� ��׾��ޠ��7�V�)iɽ�*<eɽ�*<e�Bk��٩f��S�H���0��x�1��2��ɽ�*<e'$��R��e�����kV�'$��R��e�����kV�f�{��t��;��f#Y���L-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�)V ٥�Dk����b����31�4�Ga�Sg�&q�-�+7^;]�r4�}6�X$d3�Sb���6�$%I,�R�.�c�؀7nB���I+}-mp1�kiO���l(ZQj)a#/�����ДVkr���>i4[�Xၓ�|��6C��K��f�b����|6f�aA��<y���$�~�w	�hF��z�^ƽK��,YD�^;]�r4�cú�=�A����/�1� ��%�2c��8�Y�Y��f�C����$ ��,K�"c��Y��q2q�R�s}�u�x��R.�R�����[vㆾ y�w��s��"�w�].��B9����>i4[�����) mgT*��+|��H�m�+\�����V��S���,8 �	Эr}�f�(x��4��#De(I�t)��YZ͆ˎ����~��l�h�/��_c�׈�}�y��y���dn'y&�*��5S���j{����̪j?WO!7ku�*l�<�MՓL>��RF�st�_��{�dĕ����'f%�=�5�7�O;CgE�����PH����ֺ�^-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��m 	����3���"`2:ގj����X��>%����`m{��v].p�d���ؒ�T�����
���8&5Z��?��S����{�oM���4�8v�u>) ���Y=�N����p���5��I�A�����G���R�ʹXr�=�H�m(o3����p��ɽ�*<e+teM�i��>��g�O��̱Z︷���̵oc^ɽ�*<e8�1���E�۠���s°���&GF�_x�'���ߔG�=��ɽ�*<e�Jv!U�����p�1K��9��q��N�#�VH���A�Y��gu:׈S�yg��VD��Y�tѥE��䅓�g � ���N�cv�����ۨ��wɽ�*<e����q�E������rɰ���k���,(nɽ�*<e��}Gδ�-�M`.�⽛$'a<��X�|�ɽ�*<eɽ�*<e�+\=G9I�|9��J���Mu�/�B2�:J�ɽ�*<e�&�|�D��Uo����3�\�H
̈.��A�?O�̛k�)G�'YV�yɽ�*<e�v��,��ɽ�*<e9�ݞR��=�j�8]������/��²�/��<�Q�E3#:%� 2]~����)m�L�"۠����GB���G(��[���k�Ķ*�D��|F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�YZ͆ˎ����F�7O��\�'���Ix@A`x����,9���S\��1��S���vT-ͬC�.�B&�M���F7�˦c��Cp ���t��l�4�۟�?�~r�=b)?��rB&�
�#2��;F'�Ka&��y��L��`�j�D��O[$ȫ�$m4�կ�ykp��uQih�]y��:���T:� �xs|�,TR�U����Px�YZ͆ˎ���� ����F�_ó����M�αR3շ7��L�fj��P��N×,3a[�S�nz��#�@^\�����F��2*3+^�/��p�i���1:4���-��kT	�W����ey_6�%v�	v�M�=����2��\�q
|�?���">�iL�B�m4�b�+����	qV!����Mη�D�����Ҍ�>���&5̊ _�q3y֬Ȯ�A�.I�F��y("��; xR�7�`U��ҫ�$;@ha�K�):\�H<xm�~�oB�!��r�T����m�D{�R;\�����?Ԡ�}�g���W���3�E)-_�:���u�4])�!a�+	2u�K�4�,|,:�VrW��Z�'%7���&�Mame+��Dy���9�tIJeg��7HDF�>5E���H�g�K��>��E��
�CK���"Uy��\u�� 3�J٣���6�iД�i%+gFڵ,�*ee�w��<ΞX��������F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)XO@����h[#�hV��� �L�ۄ�a$XZ�_1����m{��v].c��8.�(>Ոu����ɽ�*<e�"Uy��\�V�W�v#@CH5x�`{ѕ5��l)Ȟ 胨RJПE�[5ɽ�*<e��
���UcjoAh�q�`V�f�Bɽ�*<eɽ�*<eRu�o�V���׷@q�ɽ�*<eɽ�*<e��5c��ɽ�*<e�_F��x�I[V��k�T<z8�Ӯ`���Xu�}�_�^�&������ɽ�*<e��
���}�&�����L��m^ھi��͗
ɽ�*<eɽ�*<e��V�uA�v�x�[�Zk��W�3�clɽ�*<eɽ�*<e �.�Qq�*����p��ɽ�*<eɽ�*<e��F��,[	?dҴ�Qm��DH`�fBɽ�*<e��8t������p����8t������p�����Ɔ��"���{��߂]0;�G�	�M��)����n��d��)%��b0��a/v�sݏ����p��O�
�����GbY�%�JПE�[5ɽ�*<e�� ���{k�d�sk3Q�k.wRG�`�����p����8t����Yr5�ŕI�(^�W8 �+N�����p��ɽ�*<e��6�+v��7���`V�f�Bɽ�*<eɽ�*<eh�&U���VDL��Lɽ�*<eɽ�*<e�� ���{k�d�sk3Q�5�F`*h�� ���A�Y��gɽ�*<e����,�4ɽ�*<e�ŕI�(^�H��cx���[[Ф�����Y/#,-m�ʋxYɽ�*<e8�1���E�1�#;�6�I[⎛���b�2��B���'c@��ɽ�*<ef�{��t�'$��R��e�_o��u��1��0Q���'�}�ٔ^qt������Q�<X�3Ѧ����YuI��Q(�>��x E�3Uo����3�>|
ϒ���t�a^��mK�,]�����v��j���!bU����T�� �d!p*�~��Ϻ��Uk��+�`�C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S��W=�u�TS�:���"�˘+�)�����Ah��X�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�T�N�:Y�?���g�HpK�FB��$�A��-8��<%`�.�CD.i�>J���  ��u��ɽ�*<e��x�h
�ڝ�1�V	�	n$�n��#�c���E7`\s[C
�V[��(�[�v��4��mZn�p�qh�A�]�"(�9%O��>=3Y��
:��{g(��Î�HXt6��y��4��<*�o�lD��
���kG��z'9՗v�r-c� /L��;�R-zo���@����%���7䄲�) �ZI��������p�������Q�.��G����{�b���.����|���
�ڝ�1�V�\,��j����s�)��y����H���5��I�A�����G���R�ʹXr�	e���)Cm��Fo�ll�Z)^��_����� �
���UcjoAh�q�`V�f�Bɽ�*<e"7�!ne*5����m���8�!�|ɽ�*<e2�eme&-��'�g�����p����8t������p���_F��x�J��E|�m;ɽ�*<eɽ�*<eClϏ,8O�:�D�^��z�0�+�yɽ�*<evS+ё@{���W?t�<�Q�E3#:%� 2]ɽ�*<e����,�4u:׈S�y��5q�Ё"L�"۠����GB���믏]Ep����ܖl-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�)V ٥�Dk/���F�C�.�B&�S�E�}WM,��Y�\��?�n�t����D�˯aïd�,�obi��a}�g����;������0W^��VM1�YZ͆ˎ��10���=EFh�X}���q��E�9{$-�o�#I���Y�����?�%�>J�5��v��'h����F����j��/&)�P�Z��1��#YZ͆ˎ��10���=J��Ö�>��oln/�:3�7P�z���X����8��E�3\ǖ��HG�9Y��\���ɓ����gA�u�(��*����U����VqV�nE�x8�U=�z[����9S�d�D��xQ��`
T�(.�5b#���C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S�ɽ�*<e����q�E���蟣��B�3/���P1޸���$Q����x���]L�Eɽ�*<e���U�8�sl�Z)^��_������ɽ�*<e�|�NH_�!w510KR�����8�!�|ɽ�*<e��5c��ɽ�*<e}�tؤ�l�k���,(nɽ�*<e��}Gδ�-��Ⱥ�;lΝ�/�+;k���,(nɽ�*<eɽ�*<e����X-�9�����3�ɽ�*<eɽ�*<e���B�&�%��W�W���Iy�ɽ�*<eɽ�*<e���S��hōG�JПE�[5ɽ�*<eɽ�*<e��
���oJ�حv�N�{���#ɽ�*<eɽ�*<eɽ�*<e��yt��s_�+�:1�����[[Ф�����4��tɽ�*<eɽ�*<e�_F��x�gƧ)����ɽ�*<eɽ�*<e�� ���{k.�]�%���׷@q�ɽ�*<eɽ�*<eT��%z��.U�[�x�ɽ�*<eP�7ٝGy�ɽ�*<eP�7ٝGy�ɽ�*<e9�ݞR��=O�
����&0���xܽ��mK�գ֪ ���N@�Ƌ=��eɽ�*<e'4M���//�%
q�sڝ�o� }�uKO��m2T ��c%�`V�f�Bɽ�*<e����@�������N�ޛfe�^C�ɽ�*<eɽ�*<e"������3ɨ��U6����+H�:���8�!�|ɽ�*<eP�7ٝGy�ɽ�*<eɽ�*<e���g�q\A얺��Bɽ�*<eɽ�*<e����X-�9N�޷bPXC3���c{ɽ�*<e�.U�[�x�ɽ�*<eɽ�*<e"������3ɨ��U6����+H�:���8�!�|ɽ�*<eɽ�*<e��}Gδ�-���\�6ɽ�*<eɽ�*<eɽ�*<e���B�V`��J,Y�F��å��[[Ф�f\���Mw�w�Eɽ�*<e'$��R��e�����kV�ɽ�*<ef�{��t�ɽ�*<ef�{��t�ɽ�*<e�+�r��y��ל
ϙ� ��G4F6[Í�A��.`ܲ�V��-1Ø5i0(���nFd>��)}X�9/�a�,��mq�s��ɽ�*<e�"Uy��\�V�W�v#@�|�0�']_�@[��]�|tֿk���,(nɽ�*<e��}Gδ�-��$Q����x���]L�Eɽ�*<eɽ�*<e��yt��s_�{��L�w��NSad��ɽ�*<eH<��T�ɽ�*<eɽ�*<e���g�q\��/�žCɽ�*<e����@��G����R_�ś��{�`V�f�Bɽ�*<eɽ�*<e����@��G����R_ھi��͗
ɽ�*<eɽ�*<e�� ���{k��#W��A�����Z(�lD>`:�$V �0�ɽ�*<eɽ�*<e �.�Qq�*{8[v�
��,�fM�ɽ�*<eɽ�*<e8�1���E�`���Xu�(9۪�c���#W��͔`�gG��Yr5ɽ�*<eu:׈S�y|��5�L/%ɽ�*<e����,�4ɽ�*<e����,�4u:׈S�y�ԣ	HP�7ٝGy����2t����X��X��0C���>MX�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�T�N�:Y�?���]�^��nɖ8�m��I5�.ɹS������b�Q���5>�V��^��G�7�����:�w9���=ެVo��:���ٛA��n×,3a[y�^�Foa���b# </�űё�L@�Y�N�����ﹷ(�����ͬM�Ռy�6��h����s�
%$����'!]r&&���|"ÝW�![��Z���t�Q�F���:=%)8�82
��t��jj�gj���'9e��w,�v�
u��'R�V�*�/rXT�qP9���S�i�s��\{Y��ˀ^�Ƶ�0p&�I�ӣ|��X��˶\Ȱk.�a]�͋���[������*f�BbL&���W�u���zC�d6����
5���&{���D#�y�ҐX��w
�i]�q�6��V��oz�mșZ&<�{nvC͎A�Kf�͢��� 2��m������`�_	댇���zQ���A�0:��}�&�gO5����|6f�aA�;^�J#�EN��rE��R���)��ffs�mU�FL=�&�K8O3��H�+�6S�2�r8�Sp1�wZ�-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��m 	����3���"`2:ގj����X��>%����`m{��v].���� ��~J�LT?�H���{���zЕ&��|JПE�[5ɽ�*<e�<�l^.$G���O�{r�l�F�7�ɽ�*<ey�?E{Я�;����t���I��z��Yr5��
���#�Â{�켞�������ޛfe�^C�ɽ�*<eɽ�*<e����A�F�%�U�.�N4�:���[ɽ�*<eɽ�*<e�0vsp����%��У�²�/�	jG{{�hھi��͗
ɽ�*<e�ngF��U e1#��T��T������p����8t������p���)�w׽�ɽ�*<eX�7A?��8Xy^��2y'��/�+;k���,(nɽ�*<e��}Gδ�-�����]�q����ɽ�*<eɽ�*<e\��hߡ�8|�t*lC6t���y�Pɽ�*<e�_F��x�M�9l�v6�r��5	]�O��7��br�Z��Ϯ�&�6S�2�r8����K����(���@33�����ɽ�*<eɽ�*<e\��hߡ�8|�t*lC60H��r�dZ�ל
ϙ� ɽ�*<e$ÞXu5�
�ڝ�1�V	�	n$�n��@��e�[1��G�T;��*E��e��bUAZɽ�*<eɽ�*<e��讛 ��a�h~0H��r�dZɽ�*<e���Ɔ��"ɽ�*<eX�7A?��8���9]�(�?V82��������tn�c�{
$k���,(nɽ�*<e��}Gδ�-v�?��Ѓ�]��1,�.��G���ʫS��LI�ɽ�*<e�\�e�=l�^a�M�#����7�quA�Y��gu:׈S�y|��5�L/%����,�4�.U�[�x����h3��.
�_F��D��k��-�)>˜y/;�)%��b0��a/v�sݏ����p��O�
�����GbY�%�JПE�[5ɽ�*<e��.'�b�kz!���>�A�Y��gɽ�*<e��G3�{u5�E��-ɽ�*<e����,�4ɽ�*<e�����n�0�0��V$Pɽ�*<e��.'�b�k�4�4)�mݵ^a�M�#�x����&��ɽ�*<e$-t�O�ǱY��3M�ť��N��ɽ�*<ef�{��t�'$��R��e�_o��u����<��ݭd��PtD���K>3���[1�_V�-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�)V ٥�DkXĐˀ���]�񋂦\�m��I5�.ɹS������b�Q�/������\t=�jk{�H���Ӌ�D����G�rR~�d�e-LƵ�0p&�YZ͆ˎ�b���=���4])�!��l��%�ɂ��� !4ʊ����F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)XkwO�&뿃Ir=Xl���`V�f�Bɽ�*<e$-t�O�m/i���wnV`��J�nQE`o�ɽ�*<e������M/U�o,����F�׫����p������n��rF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�M��X�{���VJUT���kpo�%T���YW�¤h����T4QZ+ZF��)��ެ×,3a[ɽ�*<e��ZG�p4�0�x��kJ����\7%���ܖɽ�*<e�����F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)Xɽ�*<eAO�Ưu$8��>�k�Ց5�^Vɽ�*<e$-t�O�{��1�;�AXB� `g����m�����p��� 7maH���v^���q)
��aTwi �H ܷD�҄ɽ�*<e�����F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)Xɽ�*<ec=y��HzЏJ.�[�~ܪ�o(�D����33�W#�Y�R"�
}�F|G���[����!��,4���?w�[-�$%��=�3�r/��vO�����@P�2pa˲ ��H��5Ѷ�$�`�ɽ�*<eIQ����G����,���+8����y&��y~h� P����G��!��)�+��;O�ɽ�*<e\E9;�J�+�W��fx����k��xV�"��tu�e+=ɽ�*<e���HGɽ�*<e�n�0:�W
��Y&@�х�Ɉ�Q7�@Q�T�K�;�/Ͳ��{����ǥ�'�t�Bɽ�*<e3��$S���Ʒ�Y�J�g���]�q[��Ur�JF*]ŉBV��13����G  o�>ɽ�*<e�����F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)Xɽ�*<e�Z��
�rc�\����J��4g�1l�XiI�����p��ɽ�*<e- >��-}:%W��9�AXB� `�P0&�ഥ[��L�)ɽ�*<eO�
����ÚTU�ߦ�AXB� `�x[���K&
��,�fM�ɽ�*<e����@���ݝ{w,��2�0���X����� ���A�Y��gu:׈S�y|��5�L/%�
�9����f�{��t��;��f#Y���L-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�)V ٥�Dk��Mg���_����\�
��)(^;]�r4)Ӈ���z��R�{�nͧ�,���	����#S�q?�a�|6f�aA�YZ͆ˎ�g����ږ,(��ј�>�]���e�}��M�õǈa{����
Z:R�kțYZ͆ˎ�91��?��n%���H=��}�fSd�t�攮]Em�}1y5�)B��w�Rl��`�������) mgT*��DL@��u;��h�Hɷ���%`�P6��5��\ �xNC1��J�[[=�@p�r�/�Yh!f�'�NyR�G�b���w{: �K�A�v��$�i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q�ݺ����Q��F�W����m���ZB����?5��������v^�W�D6�f,׫����� ��13��91��?���"��m�
9���g�H��2��h"	H /�)�ֵb+�@���GB���믏]Ep���En�M'4M���//�%
q�sڝ�o� }�uKO��m2T ��c%�`V�f�Bɽ�*<e3ƹq�nNsd�p�{nɽ�*<e�&�|�D��Uo����3�>|
ϒ����E��o��ɽ�*<ewp���	JПE�[5ɽ�*<e�&�|�D��Uo����3�>|
ϒ���d�N(���i�yZ"c�O�K�,]�����;�:��'��l��͋��-�i:�-ɽ�*<e��
���hōG�JПE�[5ɽ�*<eɽ�*<e,�H��B".�����"�[�e�T�Ba&㓸�r5S v�*�ɽ�*<eɽ�*<e�̃n	��]�0������y�^5)��ɽ�*<eɽ�*<e1��0ɽ�*<e1��0P�7ٝGy�T��%zؕ��g�q\i�>J���6�/�ٚ(-U877�P�����h3���*�Ӈ�k���,(nɽ�*<e���YuI�$@�՛׫�*>v�G}?t�2�u��7�(b=�L��0���B��8t���ɖY׎��ɖY׎��g�H0C���>MX�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�T�N�:Y�?6�p��tjvN�yq�̭�e�Ǎ���'�K��l� mgT*�ɷ�U��8P,���\�� ��
��h�=)" ���,av���q+�aK��C| i!���l(ZQ���a�ٍx]���e�}��2�GJN����#�V�Y�y����u���vM��.9o�N�
}�X��|q�I1��*�7�����y�_Q�v��-��{nvC͎�$��!�Ng�?�9�QgH���ڄTL��~k�h�X��v���u��AP��Jc0��c�U��L�,|,:�K�235�gƦ|�c*����`��T���<�^ݻVHӽ&�����J�8���+�ތ�w���A,�w�&��G�/�����
+�6��V�vr)bz6)�X����FU���滲?8g9��;�90�DMy�w����Eڭ�{�������U#���S�5��6��u�RQh��!؈��p4��j��ڊk��Q�ryŇi�}�WC��>�����~Ð)�q�Kf�4��!��ێ�u��O��s���^��=-$Bf��[�ǧ�-4��@R�Oo,�Q�ryŇ����N���R��-�7d{�M3�s ����eP+�"�y���$`�EZ�wv�5��6��u$0��a!]N7�NK@����ZC;��^;]�r4DG��#�WA���`~����M<l28�M`�EZ�wv)#p?m-���������&��()�^k�ʱ�����u�|R��1�wF��&`��U�s/�%�@p?�&KrzJ;��U�Q�p�r�VJCW�m�L�G7�
�b+8�ԫ9�P)�`��,ch�Y,�"'5@B�A=z10,$,d�"��!�����Z<P��+�}��p��)�-� mgT*�ɷ�U��8P,���\����S�랫���Q*H��a	܅�?ru��mN�6Ǳ� W�@?=��!̶P�g%oY.3�)7Yi�8E�����8��~)5_̼�8���Au�i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q��Xƻ�2��MJ��~B*�h;��{fD��l�~��C3���c{�
Q�wP�%�������h3��.
�_F��D��k��-�)>˜y/;�)%��b0��a/v�sݏ����p��O�
�����GbY�%�JПE�[5ɽ�*<e���&B��2���m�9'�ژ`Nɽ�*<eɽ�*<e,��2�0���X�Q�NA�Y��gu:׈S�y|��5�L/%�ŕI�(^�W8 �+N�����p��ɽ�*<e ٘T{Q���v^�3�^�&���`V�f�Bɽ�*<eɽ�*<e��)����( �ͻdf/���)�6Cr��H�ƻ��on�!�Cr�4�n��mf�yɽ�*<eɽ�*<e�����߿�wL?z��G���`���t�x�x�1��2��ɽ�*<e'$��R��e�����kV�'$��R��e�����kV�f�{��t�f�{��t�wp���	��GB���믏]Ep�1<L�_ӔkwO�&뿃Ir=Xl���`V�f�Bɽ�*<e��)�������IY^����G�����-��<�WV
v��ɽ�*<e@.F�rqD�K{�utܼ�ݝ{w,��2�0����Z�!���8t���ɖY׎��ɖY׎��g�H0C���>MX�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�T�N�:Y�?ے56�{Dz����/�{nvC͎z�# �X>̡�wg?z3�t���F�9%`�ՙ9(@���&?�,��SռG  o�>H��gR���![��Z��O��tg�d���CC���+&G��Ц�L��_��Nm�j�WS�%��o��qI�K�����HG$��ƥz����5N~���;��0_�e��6�I[�O�+bjJ>&^�7�T�+ �Q�p�r�V=Ml&4��؅�(�x>Ԫ��@�)�TT��z9ტ^.|�M7N�
}�X�O0��ؾ�?'���J��ԯy��q��,�E�09���S7R�ύ"'Т���N����ԓ���i�,av�\��Y��+�Nu�&�b6M��->D�j��@�[|A����]n�M��zr.7N(OOp?�D�,�L�N+�����p�x�)�T?,�Q��L Ƶ���>�~�{�ν�&�۾��x� K��������N��5# �9�x8�U=�z�`�w$�P�-�<���{nvC͎���4zm��
ɷ'�����wꤹg?����BqOS%iv��8A��/\�V�T�%���YZ͆ˎ�!h�|�Q��2/NLa.���T8�~�6fY�l�U@O��A���(I�[L��x����,�q��s'�����b:iU�*�D��|F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��ob���O���-��њ}6�P�;�$�L>d�C3���c{�
Q�w?�-�PgE%�?�Vl��n;�e(<�KB0��Y�����p�������Q���jm��+�7��-�ߔG�=��~N�*�xʓ\[ ��J�CԶ�y6�.苢��w�ɽ�*<e�]'E���i��ѪM��u~�y‡���_����EG�r�[0�"�����޶(:�J4�2�|ɽ�*<e-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��l��q�,4���?w ��dn�ݫ)��(B86b�o�9��~T�u2��
y�F!R�0t�<Pk(���	؅�(�x>q�i�K��,4���?w���3%��"t#H�a+��*넜Th�K�am@��M�%�7"��|� -��(�'�~�uE�n�ɽ�*<ej	�%w\��ٞ1�{wz�i��F۶dlpr��������3%�"d�'5,ms�:��%\��Dy���9ɽ�*<e�5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^ɽ�*<e'4M���//�%
q�sڝ�o� }�uKO��m2T ��c%�`V�f�Bɽ�*<e����@�������N�ޛfe�^C�ɽ�*<eɽ�*<eR:�sg�
r��O�u�alZ	�%�m\6�"�NSad��ɽ�*<e�Y�tѥE��䅓�g ������ɽ�*<e��
�����8�	�`V�f�Bɽ�*<eɽ�*<e:j���+�$κp�*l|�on_�4 F0�FJ�Ⱑ{��~S*H���gZ�$M7���m���rɳ'ԙɽ�*<eɽ�*<e��}Gδ�-���q�ޤ�/�ۣ��ɽ�*<eɽ�*<eɽ�*<eR:�sg�
r��O�u�alZ	�%�m\6�"�NSad��ɽ�*<e'$��R��e�����kV�ɽ�*<ef�{��t�ɽ�*<e�v��,��ɽ�*<e���h3��.
�_F��D��k��-�)>˜y/;�)%��b0��a/v�sݏ����p��ɽ�*<e���U�8�sl�Z)^��_������ɽ�*<eC!m�C��� oISo����&��ؓ���8�!�|ɽ�*<eT��%z�s����+�P:�힗���}*.�JПE�[5ɽ�*<eɽ�*<eE�Ƹ]��'T�e~^��X5�(i�Ad��Q#N����$κp�*l|�on_��z�=�#�����p��ɽ�*<eO�
����E�R���t)ɽ�*<eɽ�*<eO@��������L3n�L��K�H֕{]�'T�e~^$��[�3�2r��O�u�alZ	��Y����0H��r�dZɽ�*<e��8t�֨��S��g�����xF�I�����ޛfe�^C�ɽ�*<eɽ�*<e�r�_`�m��ZL��!_>��d`C�����L34��?,4O���-�8wɽ�*<e'$��R��eL�"۠��Ű�����lK��H2�Sҝ�γ�������ɽ�*<eC!m�C��� oISo����&��ؓ���>j!aލ�\g��q��D�����p��ɽ�*<e�+�r��y�ɽ�*<e���Ɔ��"u:׈S�y��L��Ԝ��XS�<)�	ɽ�*<e'4M���//�%
q�sڝ�o� }�uKO��m2T ��c%�`V�f�Bɽ�*<e����@�������N�@r���28ɽ�*<eO@��������L3n�L��K���g���ɽ�*<e�_F��x�z�8ft{hc7B��ne�;����m�$V}��sھi��͗
ɽ�*<eC!m�C��� oISo����&��ؓ�@�I�����ѪM���ѬF�`ɽ�*<eɽ�*<e���g�q\��/�žCɽ�*<eO@��������L3�4}�?�g1� ^j�!ɘ�j)#��^5)��ɽ�*<eɽ�*<e�r�_`�m��ZL��!_T.�k��q��� E�g�b���rm��JVڜ_�uylZ���U��,��=�.{@<}ɽ�*<eP�7ٝGy�ɽ�*<eP�7ٝGy�����p�����Ɔ��"���{���zЕ&��|JПE�[5ɽ�*<eDǭ�\@z��A�y�����L3�O%�o2�����p��O�
�����>\�^b���LD�r?����.��Fɽ�*<eP0;g5e�:����\�� �H֕{]�'T�e~^H�6�3j��9�<Ѻ�Q�/
�#�����͕p+�2{��8t���ɖY׎�Һ��F�Y��f�2�
Q�w��$�y�����p���"Uy��\=�B��YX����p��P0;g5e�:����\�� ���g�����8t��~����)m���d�
��	D�ܣ{UW,M�d|�闈�g�HpK�FB��1�@ͫ��tiʷ����d��PtD���K>3��Će���������Q��Y!���n ��S��v>-V>�q4a�Xy�����^�}]���Iv4�4�x����(���_0( �L���y���(�nf������Q��Y!���n ��S��v>�p�G�����/ַƭ7X>��Y�8�����Cz��(I����Ph=��t��ob˒���X�i�>J���!��KR�/�j�8]��l��8��Xȡ�m�sE��@�F;}&���f�+H:lG�1G��0�'.f	&�`4�(X�/P�7ٝGy� �.�Qq�**3ZC�q�8G�X�ohX�Wk�k�s����Od���g�������0b��*��-`�C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S�4��!����:39���!� �=k��iB���u�9��J�@����z��?�3.�+�^;]�r4XĐˀ����2`���\��?�n����_I0(�S���҆�+r�GT�t�3���������ϖ���8ɾey$��]���f-dub���6"j���-(_ mgT*�ɷ�U��8P#=	
�/,�	��J�x��1و�d�F�m �
��RqR~��&Z,���'3{:^/a��f���3�]6��fJ���Y�N����p��J��d�5�Xo��e-����<�)�hlI-�-�m�
| ����&�G��7*�u>�͑��jC��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S�T`�(O��y�~�k��v���*�1��I�ۿww�Zou�_6�� ���NǚΏ�h}��PjH�U���K#�	a��}G�%4{�n�*3ZC�q�"�9u��夣�P1޸��tf�� r']_�@[��]�|tֿk���,(n��
���UcjoAh�q�`V�f�Bɽ�*<e���=c�hzc�&�c���]�֙$Dj��e�
���A"¥R>��S�i��G�-*�5fxɽ�*<e�6�/��T�Xȡ�m]�֙$D�x48802�����p��:j���+�5�N���\#���Dx뿠Z�]���8�!�|ɽ�*<e�7�=b�>����b�!�Z���E��o��ɽ�*<ev��P-��I��P�6;7}49�iv (Ă����9A�Y��gɽ�*<e�AgE	�2�ɽ�*<evE{��l��O�pٺe�ɽ�*<e����,�4ɽ�*<e���g�q\��/�žCɽ�*<e?Bp�Hy:͗4��]Q��x���]L�Eɽ�*<ev��P-��I��P�6;7}�]y\��p_xZ��C�ɽ�*<e��}Gδ�-�� �v��V�,�J�ھi��͗
ɽ�*<e9���(7�l���SIyk��X8�_��@�Y��l��͋c#ܱ�Q����p��ɽ�*<e���S���w�)�F��ƭĲ`��ּ��r=��ɽ�*<eɽ�*<e�F�.��I��'�Bp٘���%5�N���\#���D�ǋI�d��ɽ�*<e'$��R��eo�
�0�C��� �v��T ��(Cھi��͗
ɽ�*<e9���(7�l���SI~�ȰG������ƣ1�QW+�_��������s=���Ԯ�2rɽ�*<e�ŕI�(^�F��Ư@ZP���t�o��$�֩�R����p��ɽ�*<ev��P-��I��P�6;7}<�-v�;������6Zg��7V���34�/kܸ1�ɽ�*<e �.�Qq�*?Bp�Hy:ͱ��
���2�><��P%ɽ�*<eɽ�*<e���CW_s�8;7v����<��ܰk'��[���!���;�Uj�[eT�'T�e~^]A#��]�ɽ�*<e�+�r��y�ɽ�*<eSE⫄ 2}�f�}��g��e�?�ֻk���,(nɽ�*<e�����Y�9ݹE�=5�4H�x���-�poR��ɽ�*<eɽ�*<e�*E�����H�vE{��l�-T��Fy�H��n�$�����sɽ�*<ewp���	�g�k�q2��4�>I�in<����ޛfe�^C�ɽ�*<eɽ�*<e�J6���~�I��L�'���Vi��z�	LR��!&���S+G��0���A�Y��gɽ�*<e��G�H�B͜%*��ىCL��8�H��n�$�+��/5�(��CP_�Sɽ�*<eP�7ٝGy�ɽ�*<e'$��R��e�4�g T?ZP���t�o�JC#0�-1V�oz�A�ɽ�*<eɽ�*<e	H_0��pO0MGa���Vi��zQ�_����i���!�)�'hs_��j����p��ɽ�*<e�S�Ї1�l�� �v��T ��(C�c���|4ɽ�*<eɽ�*<e\e*��dX���X,�{�����Iܲͧ�0�w`^|��]`��@��9�N�ɽ�*<e��8t���)�w׽�ɽ�*<e1��0����,�4����,�4SE⫄ 2}ɍo��T�3uUrD�|!�d�٠�;��������Z){Q����4o_��8v�u>) !�-;!F��z��� ��}��PjH�U���K#�	a��}G�%4{�n�*3ZC�q�"�9u��夣�P1޸��tf�� r']_�@[��]�|tֿk���,(n��
���UcjoAh�q�`V�f�Bɽ�*<e���=c�hzc�&�c���]�֙$Dj��e�
���A"¥R>��S�i��G�-*�5fxɽ�*<e�6�/��T�Xȡ�m]�֙$D�x48802�����p��:j���+�Y��]��J��b��M&��x��F!���8�!�|u:׈S�y|��5�L/% �.�Qq�*�`V�f�Bɽ�*<e��}Gδ�-�F�.��ޛfe�^C�ɽ�*<eɽ�*<e�F�.��I��'�������wɽ�*<e����@��+�^(YS��2��4�>I����.��Fɽ�*<eɽ�*<ee�(�%O]N�kZN)ޢX���_s|�� ��!T$�����T��Z���o����p��ɽ�*<e���S���w�)�F��ƭĲ`���2�COm�ɽ�*<eɽ�*<e�F�.��I��'������DX��Wo�L�����U�ǋI�d��ɽ�*<e'$��R��eo�
�0�C��� �v���ǈ���ھi��͗
ɽ�*<e9���(7�l���SI���G'@�J� ��a���9�<Ѻ�:����~��9&ٲ��B�f���Eɽ�*<eP�7ٝGy�ɽ�*<e�_F��x�Β��\x;�g���U�`V�f�Bɽ�*<e��
���q��P�jo,b���ݮ�{U�b
ɽ�*<eɽ�*<ey�]�Ɵ�l�~�«V���34�1U����!&���S+G��0���A�Y��gɽ�*<e���S��q��P�jo,b���ݹi��H;9ɽ�*<eɽ�*<e	H_0����Iv4�4F�Kl��TQ�_����i���!�)�'hs_��j����p��u:׈S�yNd"�O������p��f�{��t���8t���ɖY׎�Һ��F�Y��f�2�
Q�wӺ��2 �K��������q�E���蟣��B�3/���P1޸���$Q����x���]L�E����@�������N�ޛfe�^C�ɽ�*<e9���(7�l���SIT0Y|:�������p��f�{��t�ɽ�*<e���S���2-�i`��ġ�Z-�}c������ɽ�*<e�F�.��I��'�V��9�pɽ�*<e��%���ݹE�=5�4�� �����p��ɽ�*<e���CW_s�8;7v����<��ܰk'��[���!���;�Uj�[eT�'T�e~^]A#��]�u:׈S�y|��5�L/%1��01��0Q���'�}�ٔ^qt������F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)XW}��Z�5�������9�R�l������rӸC��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S�!����M��%Zt݁dD,÷���R`�ߵ���1����c��T�ž>*b���寡�×,3a[�PXi=�V���34���+�%��$;����8�ђx�b9����۔�Rۢ�����Ah��mr7��;�D�b����¾_�s�̥�`��Dp�zR=�kDX~[�=Xƻ�2��U�B��뼓\[ ��J�CԶ�y6�d��PtD���K>3��Ĭ�?Ul�gg�����Q��Y�bKJ+�]�֙$D��k�!������l��9=��n�CNK퐾I��L�'���Vi��zք �7��#M��f@q7��������Q��Y�bKJ+�\�,T��aӰ����m�0k�=�Q�p����(-xc$��,Wo�5T�q�$������M��.Wj�s�8���(�[�v��.���帨S9�R�l����*��O5�Nkl��T�T�0.�z͵�$�z��3�����������5Jv`�=�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�`��ՠ~̚*D?0�:hҙ'H.����m/�D®S�&��*3ZC�q�����wf��F�߂�h5�.P�G��Q<Kt�^tD����F�W����c���C!���K�am@�p���b�!׺����Q���P'�8O�3���f��<���>;\B��Y ��!o<lr�������d<���J�ܰ�r�j�8]����ס��|�C�Ύ�ɽ�*<eF� �M��� 2G�H�m?�Gܝ�5�n�(,�[�>i �}��Pj�$�M��=l��[o �[�s�l�2�!J91��?���n�����Z��L{M�y0��bm�B���p���b�!׺����Q�`����v��]3}7�� � "a�>|
ϒ���Ț����@�U'4b_�4G������rO�^p=�(��Î�HXM�9K�r�X{�YyB���V��NENf�`����Yd��Y�bKJ+�����Љ�.�z͵�$V���34`�d��j3mli��s;E�����Y,4���?w�v�@�ߎ43�-!c(vLP���9V�3o��t���֓ߟΟ[�.Hn�G����h3��.
�_F��D��k��-�)>˜y/;�)%��b0��a/v�sݏ����p�����U�8�sl�Z)^��_�������.C��,�M�	 {���x��F!���8�!�|t9��v�ȸI��l?��
5����.�E��-ɽ�*<e̈�!��3��������e��:}ɽ�*<e��nE�$,���]@B7ل:�����A�Y��g�.C��,�Z~�;A��>��A�����-�8wɽ�*<e���cT�B\o�q��x��G��Mc__xZ��C�C!m�C��� oISo���%����r�F�]�o[��?��x��_���O�pٺe�ɽ�*<e1��0 �.�Qq�*�`V�f�Bɽ�*<e���>j!aލ�\g��q��Y�
D�I���jV���34�<k��Z��Ad�����
Jz5�N���\#���D�@��	=ɽ�*<e��s���5����_���Ei�����ݖ�>̴�-�a�������@��8��q��[����COb��{�-ɽ�*<e{�/O�s<u[�֓h�&����l�\!����ɽ�*<es����+��3I�^����[o �[�������הq��Qy�-��C�ɽ�*<e{�/O�s<u[�֓h�&����l`��X�s�Jɽ�*<e+teM�i����T� W�Cb/g���t��@0���B���¦�Гp�!�$V}��s�x{�������p����G�H�Bq5������|4�#�ol|ٖ�H^�D�ɽ�*<e�.C��,�Z~�;A��(���� A�Y��g��
���\-U3�?�dc����ɽ�*<et9��v�ȋWk��?g�%�m\6�"��
:��{gɽ�*<eؼ��y^�ɽ�*<e��G�H�Bהq��Qy�Ԍ_��4�t���y�P'$��R��e�����kV��_F��x��V�n`ny`�2��^���Z���:�j��(�$V}��s�Šs_2>����|�i41�����p����G�H�Bq5������|4�#�ol|GY��J�hɽ�*<e��}Gδ�-|4�#�ol|��[�	�ɽ�*<e��G�H�Bהq��Qy��OA�m�%��
:��{gɽ�*<eؼ��y^�ɽ�*<e��G�H�Bהq��Qy��OA�m�%�\!����ɽ�*<e�C�~�t��&�?!x�Zp���ɽ�*<e8ʦ���GWo�5T�qc�l͘Z�C
�V[�'$��R��eU877�P��ɽ�*<e!���_|�I''o�"K{E�6��h#A�Y��gP�7ٝGy�����p��$ÞXu5�nл}Z�}��z�i��ɽ�*<e�;�꽁G��
��c�MV�H
E#LPA�Y��g �.�Qq�*+teM�i����T�$9pw��ɽ�*<e�.C��,�L<�/S@�����Sb�t���y�P��8t���&Nꊓ�H�_o��u��W� ����t&՗��PY@eq�L��*3ZC�q�"�9u��夣�P1޸��tf�� r']_�@[��]�|tֿk���,(n��}Gδ�-��$Q����x���]L�E�p\�Ì���wn3�>����g���'$��R��e+�[{�����$0@��$jA�Y��g����,�4�ŕI�(^�W8 �+N�����p��X�g-a������b�C���1�Q%�����,��t~����O�
������PRٿc�ۘ�b�����Yr5�J�@1����R�Gf.h�ZI�����ߔG�=��rL۪w�Ib����?<p
����~QkRN�ɽ�*<e���䞚�/�Q ��v֕����L~_04z�9�������4�;ք|��5�L/%��}Gδ�-o�BUzZ*;�p��0�����3�'$��R��e+�[{����@B־��_t���y�P'$��R��eo�
�0�C��%6p�}��{�ć��7�ٔ�
��c�MVH[�e��N��5����ھi��͗
�e�b�-��IzJ8U݊ ���$�rɳ'ԙP�7ٝGy�u:׈S�yg��VD������Q��*E���C��,��*E�����H���?����{�nZH[�e��N�3 �\��~�3���I�[����CObX�T@}7��ɽ�*<eɽ�*<eɽ�*<e����͔߀�@sX��r��`�V�i7	��h�ǳ�y�|�-E���!��0k�=�i �*E�@�ߔG�=��h��]L�S�/�a�hd���y��UU�8�(���V8��+ Z0V��l�����<���^�=�<_%μ�R��L�����ɖY׎�Һ��F�Y��f�2�
Q�w��[u�*3ZC�q��'B�ͣ��7�(b=�L�f�Žz ��rɳ'ԙ}��Pjr��Ja�����&e�����@z�JO�
����|θ������?�H<k8ھi��͗
}��Pj���������P�h��\!���� �.�Qq�*����p�������Q�v�?���-�JCr���];��2ن��<1Ťl5��?����_0(B,���m��5�o����M���|�5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^�w����G=�_w��VS��N��>?������q1hV����qU'CU�-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�I�-��؄Ч"��+�~�K�|����%xf�R�����p���IQ����U�@Q	��
�O����ly�[��z|�Χm��ߔG�=��	t�nQ�ɽ�*<eq)�_��C
�V[�m��p�	�_@}���^� �8+�ɽ�*<e��3���/���<�ޛfe�^C�ɽ�*<eɽ�*<e�/�����ez�,U�n[�` -A�{)����p��ɽ�*<e�b<<��4r[�r�Z1BC
�V[�'$��R��e�����kV�f�{��t���FLE+����kp�l}Rk!��^�(
P��J�2�6��	�//:����#�>��xl�(T�飳������?ʌ�of�F��i��e��}R�|��W��A��1�����k{��Ty}�zj�"��0��U��j )���.s���2D��%_�y��N�[\��NT��>n.r�P�S��И]h����,��D�se��L���Ӡ��B:l��9q؟��?��6\F�߉�}3z�s"P�A/5���{�)J�ɷ�b���Ւ�tU#�݅�Cs����myW2��KqM�qsdu��&� �r��j%g�*E�Z��(wRET�1�ZAů� ��Ö|�o�l&��H�J�9B�ˎ�U�X���!4��x�ٷ�?��Ŵt� ��R����a��'��FL�j�4F�tˎ3I��(��Hk�p�IwЈ�#oԓ`��Z���GD����4�fgHg)%�RPz
2����$_�>U�V�Q���L�˷P�B�p1����Z��U�`6�!R�4�t���!���8��`�w$�P��j�:�cb�S���mheˣ��|>X,1��>�5T�g�'y{�I��y3AL�����~ָ���}R�|��`iX��-�����I���#^2�}G+�����uP�M�z�ڽS7��v�����
����%�z�M	!��Ɋn�]#�$u�	8'x��)�)�����y�>�t�Jд��߿Kv���������0���L��J���n�+cb�p�f8��H�\=҉7�#�?hX� ]����f�y���Wt�b=�D2�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�]^�h�����֖��Ws�#ג�+��n�mr$_a���F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S� h�����\��^�9�>��vf�Vg��ˉ�|<b�m���b��l�ʶ������#m�n5�!��b��i��<�a�]����2ꀻS� �]6�6�</k�M͸8yw�T��t;!7�W�<o;Gv~YE_��R"u͸8yw�T�ԍ���z��F�0�[��������\�u�<T_�R���9yB=�u�@3�2���<N�i��@����p~rև�[����9ߍ��=U
�S����?C,4���?wʉ$�Hl��1�w��A��&�|�D��.�^<�
:�ɽ�*<e���.���5��Oh`�wo�	h�[vS+ё@[;6pד,4���?wʉ$�Hl�Y}�c�oA�
+c;���)K�&�|�D��.�^<�
:�ɽ�*<e��g]�?�g��K[%����W<:K��{v���]�P�.�F� ���	/���&B�����9���P�SA����x���,�%#B����N����OQmK��h�,�B��}C��v��B��6�����`.}]�P�.�F�f�[>���ɽ�*<e{M�y0��bm�B���^�����򢋫�N���6����=���!�2X��˃�6��Rbx(r�	A�������a���D9$5U���F�����{72L%hQQ��p��u��d��q�Ӭg��K[%���~��Wɽ�*<eƚ������=��c��v�F��7 Z��B�a�h��p���yd�8�ꜟ�An0��?�i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S����>��ɝ:������ti<8=�yQaX�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8����T%�g'N�ʆQ'�&*�]u���h 0JLE��r[��h��u��ּ�&*�]u��s�(J��jf��걙I��n�_������9�͡5o�b:W�`6S�y���R)��ML�\�ӱ#�1�C�N���+�
¡$�t/"�प V%8���:��gp��
��|A�tn|I8}��]��'fj����~6��)!�������]!�I��FV�  	�F��4��Rt��A)�^U�C�y��ֳ����ɪl�VUQ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q��=�%�>}6�֮Be�%c�^Od��X�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8����T%�g'�(�[�v��9��<����$�+��� �Q�R� 	�6����^��Zlkk@�e�Yg�Sgw4���������4;���΋�q�Qy[�^N&}f(4g���?F?
fT�,p���G�����S��c^���}��Pj�p�%Ķo�
�����������rz����/�M�exْ%e����FL��>*�������1����}<@�� �� �Q~ ;z>�T-�̨� I�iE�X��X��1A���V'�i7|2d>7ε�N�SȰJПE�[55���eߵ���D~L���Љ�U&�M�OA[T�})��1���� ;�'4M���//�%
q�sڝ�o� }�DLc�w��6]�9������L����Ę�cr�����cδ�C:Z���/�žC?�p�1�}|�͆�~9��x��F!���8�!�|]�P�.�F"�#F��8��D��R����g������&B���V��P �޸����of�E��-T��%zؕ��g�q\��/�žC��()�^����5&9�B�`�b��x[���K&��&�ѯ�QPVhf(��xɽ�*<e�4R����ɦk����sW�±�����`V�f�Bɽ�*<e3ƹq�nNs��V��q���b����/�žCɽ�*<e�H��♓Ђң.���^����tQg��E.|�%���E�g�o�9�#fS�+�)���{B���h�|.U0���-ɽ�*<e�B���3�^�&��/̺�i ���4##������8�!�|ɽ�*<e��<��ݭ�`V�f�Bɽ�*<e��
�����7���u���� Q�ˀ9Ph�(�X�_���I#�L��~A�Y��gɽ�*<e��*D�g���� Q��]�P�.�F"�#F��8��D��R����Iy�ɽ�*<e��}Gδ�-���x(�iL�q�e���tseQ,�ٰ���˫�ՅM�)���ɽ�*<eP�7ٝGy�ɽ�*<e��}Gδ�-Awo��o�>���ׂ���Z�|�[JПE�[5ɽ�*<e]�P�.�F"�#F��8��D��R����g���ɽ�*<e��!�2X��˃�6��Rb��uCdZ���8�!�|ɽ�*<e��5c��u:׈S�y|��5�L/%3��֪��(���9�r���#�c�;�·-�O���#1������gW�F���>|
ϒ��޸s8����*�Ӈ�k���,(n3�5B��������G��ȓ��G,�.m��KFJ)bz1�2�+SS��g#ցi���J�KI�{O��e�:cy���YV,:��ff;R;K���1�~�#L��<�h(�ٌ�,��(:��kJ��g�-C�����hd�Fq�,��}�@�Hv@������ ��͔��\fAu=ϝI?*��cJ+����P�5���	��o��̱Z︷ko��b�e�����Y,4���?w91��?�����������F�f�x$��ʒ ��N��u�y�%E��.���Y��tL�|6�?�S�v8q�B9�*�C
Wi/��`m�i����<i��@���t�{ï|���jƤj�*4W>2��ʡ���J�#pqA��,4���?w@�󱦧�!�2X��f�2N�2���NSad��]L���z�W�D6�fg�IGL��(�I�.L;�x[���K&���j;�����p��[����Eh�.+i�b����p��O�
�����r~���.���
�BmT�I�j��5��9��P�������=��zȝ.������a�=Շ�A�Y��g1��0�my�odK���$��>r�X�gH�1�v��,����<��ݭ�`V�f�B�(�[�v��d���gˀh���D���Uv/�sbH\B�\:�y:��MH�89$)y:�I�b{0MV ��.��>�ϋݴv�x����r�ըF~�/�"�9u��夣�P1޸��ϝ<��Uצt��y4��"���JПE�[5��}Gδ�-�HYd����ޛfe�^C�ɽ�*<e/̺�i ���4##������8�!�|���ȓ]�0�D��]�-�a�K����8�!�|���ȓ]�@�r�t�O'<���ܕ�\�E��o��ɽ�*<e{M�y0��bm�B�������Bo�ɽ�*<ee&����h�V8��+ Z�E��o����8t��}�tؤ�l�k���,(n����n��r�'�)H�]@�UTv��P� ��z�|X�,|)��ٴ���ALɽ�*<e+teM�i���^tD����F�W����ޛfe�^C�ɽ�*<e��}Gδ�-&*�]u���!�P��k���,(nɽ�*<e\��I�w������-w%x�iI'������_�˭�����K�r�G�_�)�k�-u
�1���_��լR_�̎ɽ�*<e*��ׅ����U�����������|0�)მ)�����hW��r����7��_m����2�eι?)�t�E��-ɽ�*<er�֏��9��W8 �+N�����p��ɽ�*<e.݉�!V�e<+�<ɽ�*<eɽ�*<e&*�]u��	�pzwsj�I#�L��~A�Y��gɽ�*<e��*D�g���� Q��ɽ�*<eɽ�*<e�g?k�Vtև̸B���L$?��^	&C
�V[�ɽ�*<e^�W�hg��}ebP��ɽ�*<eɽ�*<eKy�1�,��K�am@��z.�1Q���D��aɽ�*<e<�ʏG�ʎL���e�Ӕ3�'Qy�c��.�ִP���K�ȕ��wN1;�ZC^����Iy�ɽ�*<e��}Gδ�-�mv�Bӝ`?�+*_�?/�}�kN�{Գ?u�̚��`�`0�B�"���dB��5��ɽ�*<e����,�4ɽ�*<e���M���r[��hlx�f8�i1E�-AEsS
/���5�C6 "�l0j�5Q��Ie�Yg�S{����������n
������1OJ���L�����'�����p��ɽ�*<e&*�]u����K�`�E��o��ɽ�*<ef�{��t�ɽ�*<e3ƹq�nNs��V��q�6|;���E�碌��V<���ܕ�\.��+(��l#b�_ީ�͆�~9��C�'Vo.#�r�f3�!1�f��4{�S�)������9���-�A��?F?
f����,q������ɽ�*<e/̺�i �>n�n���Bkv^���NSad��'$��R��e�����kV�����@��)��(�@�ۉ��i�\91��?�����j;�����p��ɽ�*<e{M�y0��bm�B�������Bo�ɽ�*<e\Jԙ�% �G������r��D��R����g���ɽ�*<e$�s�w߿.'$��R��e�����kV��+�r��y�9�ݞR��=YB8d�J5ŹG��.^Eg��Ɲ~��,`:J2�b�Y5+a91��?���9a�������[��Ƹx���]L�E~4�R�T��Q���zţ����r�[���{>|
ϒ����p�G���}Gδ�- ��\bm'���� qXEߵW�,EW ����ᠻ��-k���,(n]�P�.�F&��N�����D��aO�
����
��F)L=<RS?i�f0�0��V$Pɽ�*<e���l��'�0�D��]�-$L�pĹ�&*�]u��s�(J��jq�e�g��&��N�����8�!�|��8t��}�tؤ�l�k���,(nɽ�*<e!s�Z�<\mT�I�je�Yg�S���s�F���F�,�mv�Bӝ`�R�K��A��V��q�,�o��v�Da�;�@<BSb���!���H��->|
ϒ����p�G�'$��R��e�����kV��+�r��y����6*�H$���/J��j
���b0.d�չ�R�`����5�o���j=s}����T�73�������q)~�(����T���$�+����0��I��:�I��'4M���//�%
q�s���]�[�JПE�[5��!�2X��,�o��v
]��v��v��,����<��ݭ#��~��h�,�B�L��%X�JПE�[5�"Uy��\�V�W�v#@CH5x�`|�L��y�w�&Z6[�ޛfe�^C���
���G�?l+����o��������n��ʌ?a;�ZC^��HF3<#y���8t��}�tؤ�l�k���,(nO�
�����^k��^[
rݎ��C�ᠻ��-k���,(nɽ�*<e�9������=��zȝ.���b��4��Cl�[�6�`EO�{jL���xD��[�jB��c��#ϒ}!�Y ,��4F&��&l�c���*O��`V�f�Bɽ�*<e���&B��M�U�帶�AB
�PcA�Y��gu:׈S�y��JAc:�n�!;�l����wN1lx�f8�i1E�-AEsS
/���5�C6 "�l0j�5Q��Ie�Yg�S{����������n
������1O�c�(��
�o��|S���|0�)�Ƶ,�<�x���]L�Eɽ�*<e�!��(�V�I��ƹ��������>۳uӟ����"PV���tN�Hɽ�*<eB��6����w��_��yB=�u�@3H�iˠj&0��(e��r���"ر�h�,�B�'^��������p����8t������p������,�4P�7ٝGy��v��,����<��ݭ���H@�.�JO'����G���R�ʹXr�I,N��o+m��Fo�lS_O��k���,(n����67d���"���JПE�[5\Jԙ�% �1�o%�����\��NSad��q�И�mJ��E|�m;ɽ�*<e+teM�i����Z��L�M`.�ޛfe�^C�ɽ�*<e��}Gδ�-&*�]u����K�`�l#b�_ީ�͆�~9��C�'Vo.#�r�f3�!1�f��4{�S�)������9���-�A��?F?
f����,q������ɽ�*<eN��p޴�Bkv^����F�vM0A�Y��gu:׈S�y��JAc:�@�9���l��?F?
f$u�7���'ǋ���Њ�o��=�|��F6_��	����A�KxJ���.#�r�f3ݟjA�?xf~�mD}�JПE�[5ɽ�*<e����n��r���[���-q�5<��ך6\5笻�<S�!!
C�8)�L��?p/B?H���sO��ң�{��Y/��,�o��v��/�žCɽ�*<eB��6���a�K��'l�X�.ɽ�*<er�֏��9��?Y/����V��q�6|;���E�?��/yzX���t��g�>~�e�Yg�S�ܴ���SKj�5Q��I��5��9�����P�ML�\�ӱ#�	�������V��qٰo����7`����'�����p��ɽ�*<etʐ�&'�y�9�p���_��#��� i8 ����[Y�ɽ�*<eB��6���a�K�N��p޴��<f
U�A�Y��gɽ�*<eB��6����~�������(��B����e��e�gܓ�ɽ�*<e�+�r��y�u:׈S�y|��5�L/%3��֪��Z_���U�P��.Z#Y���L}Rk!��^�(
P�����t����	�//:����#�>��xl�(T�飳������?ʌ�of�F��i��e��}R�|��W��A��1�����k{��Ty}�zj�"��0��U��j )���.s���2D��%_�y��N�[\��NT��>n.r�P�S��И]h����,��D�se��L���Ӡ��B:l��9q؟��?��6\F�߉�}3z�s"P�A/5���{�)J�ɷ�b���Ւ�tU#�݅�Cs����myW2��KqM�qsdu��&� �r��j%g�*E�Z��(wRET�1�ZAů� ��Ö|�o�l&��H�J�9B�ˎ�U�X���!4��x�ٷ�?��Ŵt� ��R����a��'��FL�j�4F�tˎ3I��(��Hk�p�IwЈ�#oԓ`��Z���GD����4�fgHg)%�RPz
2����$_�>U�V�Q���L�˷P�B�p1����Z��U�`6�!R�4�t���!���8��`�w$�P��j�:�cb�S���mheˣ��|>X,1��>�5T�g�'y{�I��y3AL�����~ָ���}R�|��`iX��-�����I���#^2�}G+�����uP�M�z�ڽS7��v�����
����%�z�M	!��Ɋn�]#�$u�	8'x��)�)�����y�>�t�Jд��߿Kv���������0���L��J���n�+cb�p�f8��H�\=҉7�#�?hX� ]����f�y���Wt���iAD{
���9I��K�l�!ڵ?�V�7���1ء�y����UMc��D���z�/<+6���W�:R7��n	j��nfm�B}��@w/�QL�L��L�g+���_a�}���P�O$*�ג$OJ�7��,v��Z����z%u=���a�ҡ����Sk�*;���>�v�E����>�d��xff�Z��>��(��dp��*��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8���ա8&�o�	rr��I�f�Ni�Q>���ě�T�t�g��g�����63%7�K�r�s�z�b=��K�X���8�i�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e!���<��l����p��ɽ�*<eɽ�*<eɽ�*<e�uy�_q�y�NI|	*ɽ�*<eɽ�*<eɽ�*<eƚ�������]��5ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M`.ᕕ��cW�ɽ�*<eɽ�*<eɽ�*<eW�\M�'�!��&��!Q]ɽ�*<eɽ�*<eɽ�*<e]�P�.�Fi��8��ɽ�*<eɽ�*<eɽ�*<e\Jԙ�% ����Ŀ�OÕ��cW�ɽ�*<eɽ�*<eɽ�*<e��3�jh��kE�ML�ɽ�*<eɽ�*<eɽ�*<e\Jԙ�% �>|
ϒ��ޕ��cW�ɽ�*<eɽ�*<eɽ�*<e���6*�H$Y�4j��ɽ�*<eɽ�*<eɽ�*<e��\���'���DF��t*�4��T�U���Ɔ[E9錎�_K�Y�R#l�`v�4�O�RJlJ��Ԙb�խ�=����)��Q�k��/�=�����xS�u�c�8О�%��3�V����~HɃ����2X�v;����J�m��fL�1��]��DF��tdw�V���v���S���xQ��ƛ_K�Y�����u�l� �elY %H��'P�6xg{D ��C��z����3>�.��k���-��\�/ԡ59�ψ���ɽ�*<eɽ�*<e�۹MK��WVbd90a�B�a�h�ɽ�*<eƚ�����|{5�������N���ɽ�*<eɽ�*<e�̱Z︷��,�=^���B�a�h�ɽ�*<eƚ������+�(�T	���� ��#*'#���|H�iˠj&Ȝ��X|�Y��H��H���B�a�h�ɽ�*<e]�P�.�FjfA2��\�I;���ɽ�*<eɽ�*<e����#��{b�ޅ
�B�a�h�ɽ�*<e]�P�.�F�T�2+��@���W<:Kɽ�*<eɽ�*<e[����Eh\|��fW�w?S�%H��'P�Ń3^"`@T�;�/�F*���ʸ�"|��8���V����z�I�M�W��l�I&06��C�-q���njL'Kh�&�BЃW�2�G�y��jM��&d�������v��|�V^4��1�T�t�g��D^p5��d�o�M&�졩�9*��ӵ�eO���b��W���X���ݎ����8i:���~lKd��sx��f*��_�EQфnäh)�B�b� ��	���Y�ǅ%�4Y]ӄ�]l�ת&��~�af��l�G��7�1
��\�Y���<ɽ�*<eɽ�*<e���1D�RtC�i�<f"5z���UZ������ɽ�*<e�&�|�D��,�����ט��e܅�w�TN���RKD�vQFɽ�*<eɽ�*<e���x���,���Z�c�W<F�y���ɽ�*<eɽ�*<e��!�2X��)�<�L���P銆���d�A|�I4�����Zɽ�*<eɽ�*<e�B�`v��O�. �������Zɽ�*<eɽ�*<e��l�G����eX�(�4�2��R�ɽ�*<eɽ�*<e��)�����_�1��y�����}�8RKD�vQFɽ�*<eɽ�*<e��g]�?�y֘	w��J�ג�P���x�hd!p*�~�����3���RtC�i�<�6�e����ܾ�6�(�,������7dEp�������Q��B�`v�����
�_�;\B��Y ������L~k�m��c\N��:t�4��A�8�X��~ԫ��G���<G���N]������)�<�L���P銆���9��e�٪`��$N��"�L�L_R�ӽ#���N��U������b�ɂ�#�li��s;E&0(mC��b����ť ��Z����VI��b+���atBҷ��cJF�1��-ȃU`H��JПE�[5,�H��B".�U`H��JПE�[5���1DR�!�X~�hH�Hl���D%H��'Pɳ}���A�Y��gkRT����l�u���^5)��T��%zؕ��g�q\��/�žC#l�a7�Z�zK��t�;"&ِt�����p��Ȝ��X|�Y���F9�`BBF�RtC�i�<�"Q�%�����1DR�!�X~�h˲v �4x8�d�	����8t���ɖY׎�F��c�^�F����$~�M��h��#.�p7�c�xkh�qť ��Z����Vw������tf�� r��9v����Ŀ�O�ޛfe�^C���}Gδ�-����#�a/v�sݏ���{��vPBB.�`d�-������H���^5)�����&B����_�f(��X����%�����u��ѥ���-#�'H�sN�q�И�mJ��E|�m;���&B����_�f(��X����%Ȝ��X|�Y7�1
����Ę�c���1c����d�i�����L������p�����x���,���Z�c�.v1,C�C|�8�ʪ�)�<�L�����8��_#f�{��t��4��.~���A�z���n
�(,�"����Ҏ^0r��9��1ٚd
[z�Ţ-���f�o��� Cbv�A:C�]�ͻlU�Ô����0Yt�FVa�(D��Ѿ�%D�M�V�xҝ�yz�n���ufʇ��t�iW
��)%8��d}��K�n�ݚJ~��5BqgB�!�T9��A( �з��Ŀ�O�{i�9��+N[#���������rz�Ԥx���j>�˼��o^��D�}K��-u^4���Z�c��oW�8��T���Ė�eF���h�O1>�BɆ��q&�:����A���b��i���sX!�Wm��C��C��B�M{!�*B�qRB��G��5$A4�ż
�Uq���A�2?*�F�s�"jU�5�]�W�1���i�m�r��j������, ��T�B�wQ9%6���\���bٱ,�=Z)
�c��E;�RtC�i�<�ר�o��9y��W�)u>bٱ,�=Zg&c��
�RtC�i�<�6�e���#oʕ9� �q�\�>��1j��y�~�k��v-�rR3p�+�X�}�y�xxj��Fh�m{��v].�ߔG�=������4\��]�찴�}0��"�ԏ
��[n��[��q f�&�a�\C�Wd�䴼��Tɽ�*<e��0���zh!�SM�V�C�o~h!�SM�٦FԆ9�y����Q�R5�+ұĩc�p ��F�ud�^��Cī\h0�;/����pأ�a\8c��Z�c�ɽ�*<e�-͉������,=���ɽ�*<eWR�={z�1����#G���L�w�_�@2z���ue2�XZ��U������b�ɂ�#�J����A�_�@2z�����~e�U2>|
ϒ��ޜb�ɂ�#�J����A�_�@2z������VY���_�f(��%�ָ�ɽ�*<e���c�=�h�(����? +D�ɽ�*<e,؏���[��=�M.*�a���ɽ�*<e�}�k��� � P�t��Q��D*�Y����p�Y�q�И�mJ��E|�m;*3ZC�q��`��$N�2���m��b���K���bMs�ꁢ�lE���^/aö�Lάo�}߽j`��P�R���Awo��o�x����&������Q���l�G�䗍1��72R�!�X~�h��d-��Ǟ�n%�/]�5�o���X����f,6��Zl�e`a�2���s(�?A�Ҏ&�Ё?m�-�,�X�Ÿ�f�2_B@�~%.DI���:��t�%2�/	J��hא�܇*9�2�\c�5��u|R���GX��a��Xڟ3�8�H�d�h���� I���}�t�wI'[]
*�J���oE����:��C�$k5p!,�7ڐ9� ��h��'i沃�Z}����Hc�9�%�\T|Aů� �B�#��t�(a�����z}�E!Ͽ���!Lؒ&�bL�.��. ����lB��,zyj���0_��A�\��B�N��%졖*��j)?��(a�����@��$�G#�ӵI�0��#Ҟ�s�-I@>������BP�\_�0'���I"ʈ�W�rB�������i0aXK��2��H����D���i�6 ��Z�)a��\ `L���c��}W�R�#C,��n�Yx���|��/_��P��r�k���g��� H]K�s��K���{T��
�7`�	�6�#'	��m�:��eH��J�	��[W�DC�"�N�?�ot�'��#~D��\��KB����VL��'�s���7K�f*���b�0qK�s��D�1d�	!4wI�o P��z9����D�����e�mu���H��H�
:��p��؋9i�^��,1DԾ����\J���H�.'a:�s�c�A �Ы���VI#�1z���x�q��Ǝ�b\[��½�#��$̆���5��0^v�'-�r�D��6�^i~��b!�t�&��9W����z��\(u�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�8�v�_�m21�z��	���L�����}��]�X�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�4)�}Uh���"ﾆ��ъ��>?��j ���T�t�g��g�����6��2��-�C��uԅsb=��K�X���hs���ߔG�=��I��&6=��a��h���͌:�\�I;���ɽ�*<e�l��m	�&�|�D��.�^<�
:�ɽ�*<e�&Z6[ߕ��cW�I��&6=�(n?�����k���\����W<:K��{v���ƚ�������]��5�F��7 Z��B�a�h�ɽ�*<e�M`.ᕕ��cW�\�I;���?��Q�~�P�f2�]�m�]ף	C"Ɔ�;��t�^	�ER���-��Ę�c5����_k`ɽ�*<e�C�.��MҼ��>i�5��M���>���6�����&B��E����Ѳ����{72L%hQQ�ܑ������my�odK���R4͑aC��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�HE��޻'���n-l�4��wy f��F=�����F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�Oњ����4�P��\b;��s������с�p�%Ķo�&��_h�Lܹ"$����C}�/��cF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^]�
��R�!<ǪEu�"īǞ_��fi�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S�*����n4CmVt.���a�:�{r��Aiq��%���G�;�E�E�[}j������y������9T�,p���G������4;�
Cj`▘9�����VA�/�l<~O~���h�M͠8�H`�����o��������Bp��P�S_O��k���,(n���ȓ]��P�۫u	�ai��#��&Nꊓ�HL�"۠��JПE�[5����@���_��u���0�S��3�^�&���`V�f�Bɽ�*<eɚ���5.��<�^�e�:��@�Re<+�<�W�0�8�͆�~9Ț����@�����,k���,(nɽ�*<e���ȓ]��P�۫u	��|5a;�D�ɽ�*<eT��%zؕ��g�q\��/�žCɽ�*<e?�p�1�}|�͆�~9�E��o��ɽ�*<ef�{��t�ɽ�*<e1��0����,�4���Ɔ��"�"Uy��\=�B��YXHv@�����b:@���������� ��Mb?ߎ���)����� 3�ä0H��r�dZ~4�R�T��Q���zţW�D6�fp�,I��_�0�}�CPm�k��~QX�j�5Q��I��5��9�ə�/5�5��zX���t��4k���o��!�2X��`p��BN��D�_���Z��a���[�Bд�>*��� ���Ғ�#����Cd4-���P�.׵���Z��ɽ�*<e"�Y�n����V��q������]<��%m (�kE�ץ��,��х!;)���ȹ�z���������$�����p��ɽ�*<eu����'��mT�I�j��5��9��,��RO��V�]��<�	�x�(aE2�M.VyN�n���I�\?�YMԝ��zg�43�Nɽ�*<eɽ�*<e��a�Iw���΋���'(f9���Bӟ�nည�����Uj�0<gn]�0���e���w�\
h�["M6f��������5�JF�M�Vy�cgͼ��UQ�N��V��G���Y���C��&�-�,�X�Ÿ�f�2_B@:P��dS	nT��e�&��F]�J�������	U�֝�%��LP�b�I�hS\'��/���`b]P�L��ϰ�9_��]-͍)�,\���� I���X�%���=��dn'y&̢���N���ꗳ�)�70bxN7~/Ǧ��!Fȵa�E�UJ̘�P���W��-�\��\����WgƘc���Jt���M���bf�\c�ꗳ�)�7�;⑤���a,�"�빱x�Q<�^eg��ɂ����c_�o� x/���C $P��!zsv|MC�[��ĺ6
&���?��������Y���i{\�M�Q#�`>�P����Yy��0�	ĭ��n�W���\?�R�?3�h0)�E�Z��(w
�7`�	�6'�����<5���K�����,%GJ�k���.Ҋ[m]1��F�^v�'-Ɨ�8;�gi��{�]<�S#��B����2"��
��V������+�v��Tj0��L�m��7���dO��H�\?�4x!�i輸m�a��&�^��=3���,je6�����B�g��o&76� ���+ɾJ�Y�WX���v�	p��i���y�6]v��P|Λ#�2�[�k�tf�����0U������J�yP��}H�{_�.�@)1�7-��H�&��_�6�*�q#�L
2�������̹�"�j��;�kԐH`�Q��
I�DYZX�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��?h�Z����Up	ȶ5�~��`�TX6�]�G^�	X�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�4)�}Uh���"ﾆ��ъ��>?��j ���T�t�g��g�����6�y���Uᷘ=s{q f�&��p��Hv@�����Uj+����1�2P'L���Ę�c5����_k`ɽ�*<e>"��;a��F��7 Z��B�a�h�ɽ�*<e�.��W�Hv@�����Uj+����}NВີ��/�žC����N���6����=�wRۣB���kE�ML�5��Oh`�wo�	h�[����@���F�f���Ę�c5����_k`�'�jZ���Y�y�Na	-H���~���?-	��1XLם�A�<��V��A3��&�|�D��.�^<�
:�ɽ�*<e��g]�?�g��K[%����W<:K��{v���]�P�.�F� ���	/���&B�����9���P�SA����x���,5b]���j�����F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�ol&���rl٫�����"�iY��6���9@�5��5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8���e�̣�9Ph�(�XJ�`Ŵϫ��A)�^U��Qew5�I,ŶU��xv��J=�l�VUQ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q��=�%�>}6�֮Be�%c�^Od��X�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8����T%�g'�(�[�v������ ��eB4�������4;�H���q�Qy[�^N�h ���ki�J���-وɴq��G���n�(貨��'4M���//�%
q�sڝ�o� }�DLc�w��6]�9������L����Ę�cr�����cδ�C:Z���/�žC?�p�1�}|�͆�~9L@���T$u:׈S�y��L��Ԝ�x���]L�E��
���wш�� ���C�L	Vހӝ3\x���]L�Eɽ�*<e�ܳ�~1�p������9�W�0�8�͆�~9ޛfe�^C�ɽ�*<eɽ�*<e/̺�i ���4##������D��aɽ�*<e��<��ݭi`�iWӤ���Z�|�[JПE�[5ɽ�*<evS+ё@��V��q١$Ϡ��A�Y��gu:׈S�y|��5�L/%f�{��t���8t��0.d�չ�R�s8����*�Ӈ�k���,(n��q�Ӭ�t�u�`�0�T�2+��@,4���?w�ۅ��1���������-E���=#)ۏG0�\�0�&�i��BfeD�d����Q�蜅��d��|;�o�q���OҨmO��f�C�xi9&*�]u��é�N����Փ�44sQ�f��(��7<�S:V�	0�3���&���&B��2���mܗ�Mϩ�fj���M���z굺�U���1z�geι?)�t�+bO!!o@�uG\|D����{f��S�H��1����}<@�� �� �Q~ ;z>�T-�̨O�. ���y���S�ӗ=E��RxT� ��i�spoz�X�}��R��Z�J���F�c�q9r�T�?:�;���A��#�P:\����u)�QX^�2���@i"M6f��������5��	"	���?��o��N�1�a�g��ۓyP������1��
O?�p٫j��"�yL�x���Ys�}�q��?Xٵ��5�,����F]�J�������	UQQ*rb�5��6��uF�p�	_�P塙@:/!M_[V�I'�
n� 70^�d�e»�-0^��,�:�	S�uP�M�zK!�g٪�'�)��F�p�	_ى�#�9�$�oWU� ����L�m�C��#��;����B�	?�gwC�N�O�lK���K)��F��P������_#Ǚ��R�����'c.�	?0-� ����Jv���,����@p~�@oH��{T��qɮ����D���,%GJ�=�rW�K�v��|�5������zWG����ʙD�0@]�����>'�6�*�q�t������ϩU�R�4�t������:Wp<!���I��d�>�r=D�9�)�Ί#|�Ӏm��!Q	s>R=��@�wG�ɽ�&���[�O�VG/"���@V��"W���à\j����f���ԝh<K��}|�?�M��\%i�������E�!��o�8���RX<���O��"P)�6�m�`�� P����Y6Z����*y����,��/�&�5K}�*���ՙ��e'�������s�SŠ��z��Qd_No���?�%6=�tg���>�C_9-���\�����"*/�ٮ$C-�}Ԧ �+�[�	ݛ�&��=���y���j2�0�F�P���5c�"H��Y�ա?���c�t%�A�}����@��D �M��H!DyX�ܞ��c@[�<l:]�y��9O�}Q�g+��.�h���J�,]j�\�v�������f28�/����<{�f�%t��ts��>D j�Y�*�'s�W_7��HDč��D�"�iS{/E�́7�׈�|�.�Q>���ě�T�t�g��g�����6�=Ff�pjca���D9$b��i���sX!��-�几��p~rև>���x��Y��,��[{[T�3E��J�(g]�nȻ���O�;k��f$E5��7Z�Eߛq+k��Õ��Uɽ�*<eɽ�*<e�VJUT���H�SQv��\�$ �2dͤ	�����|d$o���vU�[��xLwq��_�c�Q�k��/�z��ʬ����<wO`r�n$��o�;\�u�<T_9��`5����[No��<wO`r�n$��o�;\�u�<T_o�:�z��}r!b&X͸8yw�T�4����^��M,�Q�.#�����{��پ�X�[{*o��^��DF��t)vD�厜1� �b�t7,4���?wP�;�� s����� �;�ū��bf�\c���G\mP���DF��t
�-P;ޛ�g�n�5�ۉ~�5��;�ū��bf�\c����01]�Ҽ�w	�I�D�J���u�|�N����>]�Ҽ�w	�I�D�J���u�| JB���T]�Ҽ�w	�I�D�J���u�|�]���M��1����{T�_0�����u�|M�iY���+]�Ҽ�w	�I�D�J���u�|�R��+�]�Ҽ�w	�I�D�J���u�|�1����"�����sʶ��6L&ꬶ�Re6R������"�����sʶ��6L&ꬶ�Re6R�����(1�;��w�)3��Z��������[��� �,�]�Ҽ�w	�I�D�J���u�|�n�[����Z�$DC����yl2����ar��Z�.�S$n�;7	b=�(|�4ƍsK�_Z��~��WRKD�vQFEŝ�h8xf���cWN7 �ϵ%[��zN�����66/�@�H[-�H���G�"�����sʶ��6L&ꬶ�R6�O�C�8J��^��@]�Ҽ�w	�I�D�J���u�|�n�[����?�^ȉ'I&�yl2����ar��Z�.�S$n�;7	b=�(|�4i\cgQK��~��WRKD�vQFEŝ�h8��l`.��N7 �ϵ%[��zN�����66/�@�H��5�
��y�\�r
�w�)3��Z��������[��� ݊&�S_V]�Ҽ�w	�I�D�J���u�|�n�[����_b���h�yl2����ar��Z�.�S$n�;7	b=�(|�4D\lU�x���~��WRKD�vQFEŝ�h8�q͜R*�{A���� �ϵ%[��zN�����66/�@�H&���D>m��K�L�V�'w�)3��Z��������[��� �мM�uS]�Ҽ�w	�I�D�J���L�X��;6V'��	w�0u�a� z_.?�PZ������M[��m6�����>�6 z_.?�Pބ,&��2M[��m6�I���8��~��WRKD�vQF�:�#;]�Ҽ�w	�I�D�J�vS+ё@[;6pד5��Oh`B�VT�́�J�@1��.8��lg��K[%���Җ LF�lT�:�����,��H�KV��iI�5��M�����x��{.�#A���Mc(J �����>��y~w�)3����Y��G���KT��&��!Q] �ϵ%[��zN�����=F9��Vac]8���}���W<:KRKD�vQFpH[��V�x����Q��ic��ݤ���S���)��i{ޝ��i�O^������(h�Ł��Җ LF�zN�����O���8��H�+o?�T�5��M�����x��{`�ܒ��eE����Ѳ�M��1����{T�_0�������_u@>R}9�ܻ���"��aa?\��E�h�,�B��,J�k�껶x�q'���M��1����{T�_0���8�1���E�F�ʔ1��J��E|B������k{sAa#�0�&V� CB�S�K
�L;��*&ꬶ�R{�F�U���zN��������؈�RKD�vQF�$�j���4�2��R����b�6�x����ޖ�zN�����!���w�2�(���"�Bz|4�ԀzN�����!���w�2�(���/��bv΀zN�����!���w�2�(����NF��q!���y��8��d��^5)��}��PjM[��m6���!�J�ڣ��g�.�k2�G�Cz�,;�T�*#�Gm���`I_{.c+O0��I���/�žC�R���.���Z��spu?�*i_�{E���D�&�T�t�g���xv�
gmǏ��m 	]�ͻlU�ËE�˵J�짩���Jp�-j�΃`�ɽ�*<eɽ�*<e��v2� +�n�/�G��|Mt"ɽ�*<e�%CX�sd���cW��b���o��ɽ�*<e[)�i�����r y!�}��0��6j���ɽ�*<e(�B)�����p���I4>���ɽ�*<e�E���s4Z��[��NVW���P���S#��\���V��oP&[<�F4h6m���(�:���[+�n�/�Gn;��w#7JK���F1�=� x�+�n�/�Gn;��w��vX���SE3�	č+�n�/�Gn;��w:��/�M��SE3�	č+�n�/�Gn;��w,�}NhG}�F1�=� x�+�n�/�Gn;��w� �g�e֟E��Q�={g����M@~��Z��ɽ�*<e- Z��(����l`.���NS���k��W�^a�2��f�������p��v\]�3OU�2�(���3/'�S���I�v�:�ߔG�=��q!���y3|wU���^5)��T��%zؕ��g�q\��/�žC�����Q���u�����P���{��(��Î�HX����~ ����;aʈ�E��(�[�v��Yγ5h7&��E@ѭYA�Y��g��x�h���.�G�6V'��(7L���������Q�n;��w ����7U;H9 K=�8��3��7�W!�s��	�J� jLⓊCf�"$�;���^/a�61�fS�7h6m���M1�?ρ�.�_C����\�3�]h}D��Y&���[��� 
r���t�*3ZC�q���x�YU$�TҘ��Sˍ�����C�6$��J�.�$3��1�����@�h}ϭ�l`.�����p�x�"�B@5�o��3����R왿��!�%�hP����)��I�L{���"��&����)��AUq�i�K��Q3��Ѓ�N䯎��eN�<v��+X��a��WD���Ɯ�h*z���c_0+�n�/�GA! �+Є��?@�����cW�ʚO�z�9�_Y�o��7�+�z��ʬ����<wO`r�nlS���=�+�n�/�Gm�K�֩XQ0)I�P�z\m���� �{����k>��E�c4����l����+��)�����u�i7|2d>7OO0��~�L���sc��O
�(D��B��;Cc�{��詐d=�Q=��V�>�}�(���X�Z�/ʛ�_�wɽ�*<e��v2� ɽ�*<ec+�V��Zɽ�*<e�%CX�sd���cW�$Ƴ¬���ɽ�*<e[)�i�����r y!+�n�/�G�  �X|Jɽ�*<e�U�J�ĕ��cW���:eA�9�W�^aǯl�SX���S#��\���V��o���V�uCM�V��L��TҘ��SIV��n;��w� �g�e�ՠ�q�1�W���P���S#��\�VV�*H��c���M��l`.�����:wd/+�n�/�G�נ�G����cWζr_�g-�������`��A��ɽ�*<e����C=�k�V��6*SD+�?M�Ȧk�v��"Rݗ]T�Żm�3'k:�@	 ��U�+��c����V�uCM5�R(�*����6���n �u�HYȦk�v��"Rݗ]T��'�09k� ͎8qRfSO�݁W/���ɽ�*<e�-�bW�����̯�B!��^7_�ŕ��cWζr_�g-�ֹ�TC�rO!��ŀy�2��Aqz����p���t�<=��ǂ'J��r9��S��*I@��d��V�pɽ�*<eċP�q�M�Q�Ğ/��ᦲc�����p�� L՚`Rp���K�`�r�fp�:�A�!�ɽ�*<eT$��t�����Q��#p��w~ɽ�*<e�����V���8t��Һ��F�YgƧ)������GB��᚝irZ������zG�J��xҦ �l�CЀ_�`��'�x 8��m�vS+ё@�Y�A.<>|
ϒ���A�Y��g��xqv�>Z]�!0��'{�5r{�]'E���i9b��no��0�(�@w�O�. ���c�0�I7�kwO�&뿃"�9u��夣�P1޸��ϝ<��Uצt��y4��"���JПE�[5ɽ�*<eBp��P�S_O��k���,(nɽ�*<e0�(�@w��X"��|����8�!�|ɽ�*<e0�(�@w��I��'�t���y�Pɽ�*<e��cE"B���BE�٫���8�!�|u:׈S�y|��5�L/% �.�Qq�*�`V�f�Bɽ�*<e�6~��T��W1�M�(��V��`��ɽ�*<e�/�(o��w_���׹�g��>��'ɽ�*<eU�8h�b�_pR/�Pɽ�*<e�W7P�%lK^���_r�P�]�ɽ�*<e�p\�Ì��H�:���"���Mɽ�*<e�wNF����2EG~�Q͎�&��!Q]ɽ�*<epH[��V�� ���	/ɽ�*<eɽ�*<e��5S�kE�ML�ɽ�*<e!ՠ��sr/�0!�$�ɽ�*<e��I�v�:����p���H>���h~�U���u:׈S�y|��5�L/%�J7�a�@������/BƷ?�yN��d3M6�3��,q��?�Vl��n���
��4P����W�Y��xlY����p��m�9���c�J�Y�l���(g����p��m�9�W���3�>Ѻ٤tF"7�!ne*5�wk+��<���t��!�]c'ҘFj�om��Q3��Ѓ�N䯎��eN�<v��+X��a��WD���Ɯ�h*z���c_0+�n�/�GA! �+Є��?@�����cW�ʚO�z�9�_Y�o��7�+�z��ʬ����<wO`r�nlS���=�+�n�/�Gm�K�֩XQ0)I�P�z\m���� �{����k>��E�c4����l����+��)�����u�i7|2d>7OO0��~�L���sc��O
�(D��B��;Cc�{��詐d=�Q=��V�>�}�(���X�Z�/ʛ�_�wɽ�*<e��v2� ɽ�*<ec+�V��Zɽ�*<e�%CX�sd���cW�$Ƴ¬���ɽ�*<e[)�i�����r y!+�n�/�G�  �X|Jɽ�*<e�U�J�ĕ��cW���:eA�9�W�^aǯl�SX���S#��\���V��o���V�uCM�V��L��TҘ��SIV��n;��w� �g�e�ՠ�q�1�W���P���S#��\�VV�*H��c���M��l`.�����:wd/+�n�/�G�נ�G����cWζr_�g-�������`��A��ɽ�*<e����C=Z�084S�����c�J�C{u�h��@����p���v��̟�}+��c��{6����hƁ�,3D>�d�+�n�/�G�n �u�HY*�W28���í�2ɽ�*<e��ٱ0+/Ð#�^���ᦲc�����p���"����#�n!@$��儙'Av�'�B����p��U��`���5 <�t-*���a��m��O^���̀2Qtf:ɽ�*<e����z	�ǂ'J��r9��S��*I@��d��V�pɽ�*<e����H�Ր3i�0X
Es�1��)Z���V�uCMN��$��	�)��¹u)^R�m�J��M�U�帶J����A�,4���?w��C�*6�	�z?���hY�����I�v�:����p������p����Q�3����BrW����Z��!�S�B���>#�{�M�ɽ�*<eb/d2��ђx� Ή�+��c� ����;�����n��;��2��:7ɽ�*<ez���y�7��,����sE��@�6��m��E�����A�Y��g���  I·���u��_a������ ����;�z�`u�t��'{�5r{,4���?w�����Q��
Yz�,c��-��|"t�H�9�� <�t-*�A�Y��gg��xK�Ҧ �l�C�8m5���	�v*��}�',0J,ͪp��b�D�D9�G�J��xҦ �l�CЀ_�`��'�ɸ8�u��}��Pjy	J�X쟋f�2N�2��0�(�@w��+�(�T	�ɽ�*<e�����Q�E%��D�&���fD���2EG~�Q��V�)i(��Î�HXV �y�l��ѥ����*�~@�gZ�T�2+��@ɽ�*<e}��Pj�j�K�Y6:�8Í�7P�\!����ɽ�*<e���I��cW�n2dꜱ+�	����p���(�[�v��Yγ5h7&��� \���NSad����?��zF�	D�ܣ{U���ɂ���6��Zl�e`�KK���o�s(�?A�Ҏ&�Ё?m�-�,�X�Ÿ�f�2_B@�~%.DI���:��t�%2�/	J��hא�܇*9�2�\c�5��u|R���GX��a��Xڟ3�8�H�d�h���� I���}�t�wI'[]
*�J���oE����:��C�$k5p!,�7ڐ9� ��h��'i沃�Z}����Hc�9�%�\T|Aů� �B�#��t�(a�����z}�E!Ͽ���!Lؒ&�bL�.��. ����lB��,zyj���0_��A�\��B�N��%졖*��j)?��(a�����@��$�G#�ӵI�0��#Ҟ�s�-I@>������BP�\_�0'���I"ʈ�W�rB�������i0aXK��2��H����D���i�6 ��Z�)a��\ `L���c��}W�R�#C,��n�Yx���|��/_��P��r�k���g��� H]K�s��K���{T��
�7`�	�6�#'	��m�:��eH��J�	��[W�DC�"�N�?�ot�'��#~D��\��KB����VL��'�s���7K�f*���b�0qK�s��D�1d�	!4wI�o P��z9����D�����e�mu���H��H�
:��p��؋9i�^��,1DԾ����\J���H�.'a:�s�c�A �Ы���VI#�1z���x�q��Ǝ�b\[��½�#��$̆���5��0^v�'-�r�D��6�^i~��b!�t�&��9W����z��\(u�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�8�v�_�m2[� �����fL��7����Y�=��/Ms)�s^#Q�&tb���F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�
�c���z��g:�Bح�xHi�����9Gt�o�iDz [[w/�QL�L���R��9E��|w�e��DZ���mq f�&�,/�z/�W�u������A>��Kji��p�ނ&�;�6���nF� �TO��ӹvji��p�ނ'�.Aw��2����άb�����O1�4{���C��DF��t���0UH�i7|2d>7P������p�(7�:Q(д�`8�1������~^-C��V����C"Ɔ�;��t�^	&2Bv�s��yl2���ɽ�*<e�G�x9��F�G��/�gj��� ��#*ɽ�*<e7��� h)��Rd�'�C"Ɔ�;��t�^	�斚IO�`�����G�~�ăC����W<:K��{v���ƚ�������]��5�F��7 Z��B�a�h�ɽ�*<e�M`.ᕕ��cW�\�I;���?��Q�~�P�f2�]���&��!Q]��~��W��	�m��yB=�u�@3�&而n��P���d�����`.}�F��7 Z��B�a�h�ɽ�*<e�(���V8��+ Z���cW�\�I;���ɽ�*<e7ӱ}�	i&�K�am@�᥀]a��?-	��1XLם�A�<��}5�:�F��7 Z��B�a�h�ɽ�*<eAwo��o�V[<Y7�0Ϣ���N���6����=���!�2X���=��c��v]�P�.�F�f�[>����p���yd��l�G�䗲Sk�𷉋5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�(���~B��ι��%J�����{!+�YXz����i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S�k��S�1�g:�.�Uݤ�}n�������x"2i7|2d>7��	׌!�J=c@�LT7~�1��k�ih��5�od���/�AyB=�u�@35�ޏ�ē[���������v����7�G2���jLB�~qO���&����>�{�?�M�U�帶�}��}���mv�Bӝ`$2���#齕�;Y5^�)�[����;t>R}9��]34/�+/�� ?��1o݁��!8�v�������a��TK�L���e��,xX�u��{v��ګՏAAz��ߘ�*JBqAktz}�{�X� $��ӣ�u�R)E�݁��!8�v������ɈW|��W������)AW�P�������x+��dԓg��V	�Pxx]:-�>T�Ǿ�*l�-@�81l���W��;�ˀC��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�HE��޻'����������L�Rh�l�VUQ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��&Ic�E̺����Q����Հ9UT�,p���"c��0Q��LX�"9uɽ�*<eɽ�*<e�&�|�D�¡�)A��I���������|v�|�ɽ�*<eɽ�*<eAiq��%�L���׫�{��ɽ�*<eɽ�*<eY�y�Na	-�kK7�4��ڬ��i(��}��Pj6���V�VۺZw/�ӽ˃�6��Rb��9s0NO�����Q�˳�Cd�2���ݝ�G5�td'�bQQ���y=����_�ņ#��偆yB=�u�@3F8o��S{�`V�f�B�ar��Z�.��U�kF��!Z�_�q�Qy[�^N&}f(4g����w�����#;�Nc���ġ��=��{�6��l�bY�t��y�������Q��81l���}�)�f�B˳�Cd�2��mb\g9-��q
C��':{�ک��"Uy��\�V�W�v#@CH5x�`|�L��y�w�&Z6[�ޛfe�^C���
���G�?l+����o��������vn^c��'�$Ϡ��A�Y��gvn^c��'��q��Y��A�Y��gvn^c��'"�h���RA�Y��gvn^c��',�o��v�E��-:j���+�Qn�g'�Z�'b)2�����g���o��Q񎑍n�≱�P?���)өֱ�E��-\Jԙ�% �f��S�H�E��-\Jԙ�% �>|
ϒ����E��o��ɽ�*<e�mv�Bӝ`vk�q嚤���8�!�|`�Uڊ%7*������W�5M�<�{���g���Y�tѥE��䅓�g [pe�2�f?��}Gδ�-Awo��o��������\Jԙ�% �>|
ϒ���b �cF���ɽ�*<e]L���z�W�D6�fg�IGL��(�I�.L;�x[���K&�ێ����ɽ�*<e91��?��u��6�������p����̺ ����U������b4�E!�:4ʛ��M��M�,W���ڀ�Jr����� �
����6���޾(lx�f8�i����)^މ��R=>pAJПE�[5ɽ�*<e����@��䛤A]��K�`_�z!�`�x���]L�Eɽ�*<eɽ�*<e�#齕�;ML�\�ӱ#=���3e�%����p��ɽ�*<e]�P�.�F��u�ǧ2�gt.�A��ɽ�*<eɽ�*<e��ɈW|��-��v�ӽ;\�6�ww��P�ߜ�v9��e�gܓ�ɽ�*<eɽ�*<e�� ?��1o6|;���E�*��,r��K�`A�Y��gɽ�*<e��
���
֮9�8WD����#�Zl���U���h�,�B�̮/�|��ޛfe�^C�ɽ�*<eɽ�*<e��ɈW|��W������3E��*�����D�ǘY�in�� �LX�"9uɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�-��V  �Y�in�� @ˀ��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�-��V  �Y�in�� �������ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�-��V  �Y�in�� ��W��������p��ɽ�*<e��8t������p��ɽ�*<er�֏��9��F��Ư@�~S��͸V/?%���-�A̮�^ �U�xJZ\Ju���/�žCɽ�*<e\Jԙ�% �f��S�H�G*�ag(DA�Y��gɽ�*<eG}�Q���еB�_3�3�,���D��aɽ�*<e��8t�֨��S���a�t2ΰo����7`�`V�f�Bɽ�*<eɽ�*<e��
����r����pQWuX.����������ɽ�*<eɽ�*<e,4���?w�'	L���3�)&(���)C:\Gt�O�����Z�:O�%��q6$��O.+��`�^/��ɽ�*<eɽ�*<eɽ�*<e��}Gδ�-�mv�Bӝ`�*]{��1l�XiI�����p��ɽ�*<eɽ�*<eɽ�*<e��}Gδ�-�mv�Bӝ`k�@���I<W�N1-�4��t��%M5�!M�u�R)E��g#!x%qgg���=0)�=E�ڎ��"�&�"Y���V�m�F@�`w�,[Tե[h27�� ���96/�>�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e<\�"��ɽ�*<eɽ�*<e���x���,8�T����[R�Ȫ��@<BSb�����qD*&a���|I1VƤiN�
�x�q\�@,��-gg���=0)�=E�ڎ��"�&���B����ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�PX���7��_m��'=n�^�ְ��yK�}Q�`Ɣ�t4���ɽ�*<eɽ�*<eɽ�*<e:j���+�L���e�ӳċ*���٨mv�Bӝ`�s�S��4���
:��{gɽ�*<eɽ�*<eɽ�*<eɽ�*<e2��Za���!���X"z�$�0-:O�%��q=���X�#�j�C:=�T�"��U�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eA�����-��v�ӽ;���0>�K�>R}9�����k%J�?��kv_�d�����p��ɽ�*<eɽ�*<eɽ�*<e:j���+��~S��͸V/?%c�ٮ:���ɽ�*<eɽ�*<eɽ�*<eɽ�*<e}�� �cۏ�d�H�*,<���ܕ�\�ՏAAz��ߘ�*JBqAktz}�{�X��g�P��J�	��H�3����u�]x)��� >���q�4����Vɽ�*<eɽ�*<eɽ�*<eɽ�*<e�y��]3%$�^�ְ��y��͊1�B�,�{�o�}��y^�=�0Ps�%B��@��6#���ߘ�*JBqAktz}�{�Xj*4 ��I@��T52�����p��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eD�*��2>n�n��]s�P?&Q5,������[�������U��,�{�o�}��y^�=��JP�$��e1��$�֜4���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�!������6|;���E�vA�=��J�	��H�3�����W���)5,������[������3�ө��A�s;�J`r7;5lrɽ�*<eɽ�*<eɽ�*<eɽ�*<e�+�r��y�ɽ�*<eɽ�*<eɽ�*<e�Y�tѥE��䅓�g ������ɽ�*<eɽ�*<eɽ�*<eB#��Ko������ GpJg@�;E��Y~�D�X������)�ܩq�8�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�ā�d䟍�������A��E��^��Xm)}Aɽ�*<eɽ�*<eɽ�*<eɽ�*<e`�Uڊ%7*������W�5M�<�{��2e��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��!�2X���I��'�l���)�8��d�H�*,<���ܕ�\�ՏAAz��ߘ�*JBqAktz}�{�X�{�,�v�n�J�	��H�3����Ҕ:b9��=�l/ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�Y�tѥE��h���y�~��\U�(D/�v��C�� ?��1o6|;���E�vA�=��J�	��H�3����:^=�A8u5,������[���&(�J�-�A�Y��gɽ�*<eɽ�*<eɽ�*<eW�h;�A��M�U�帶o������ɽ�*<eɽ�*<eɽ�*<eu:׈S�y|��5�L/%ɽ�*<eɽ�*<e�q�И�mJ��E|�m;ɽ�*<eɽ�*<eɽ�*<e��}Gδ�-�mv�Bӝ`k�@���Ii�
��T���Yr5ɽ�*<eɽ�*<eɽ�*<e��U�kF���p#n�[AK>A��kN��Yr5ɽ�*<eɽ�*<eɽ�*<e���x���,�V8�K��,�o��v^F��$'��Yr5ɽ�*<eɽ�*<eu:׈S�yu�Ƀ��M�f��S�H 鳠⃅�Y5^�)�ɽ�*<eɽ�*<eɽ�*<evn^c��',�o��vdB��5��ɽ�*<eɽ�*<e��8t������p��ɽ�*<e����,�4ɽ�*<er�֏��9���rr����&a�(j;���r)_�/�� ��/�žCɽ�*<e�H)��k�F��ɱ8\C
�V[�ɽ�*<e��!�2X���I��'�B���A�ɽ�*<eT��%z�s����+S"C�J
��3/�})�޷����wx���]L�Eɽ�*<eo��Q񎑍�\=�6���Iy�ɽ�*<e���&B��~��\U�(�gƋ@����ߔG�=��u:׈S�y��JAc:���V	�2��1���`"��Vd��)'�`V�f�Bɽ�*<eɽ�*<egR&O�)1*f&�Rk��ɽ�*<eɽ�*<e��l�G���/}�Ofgٹ�`�7.\�'$��R��eL�"۠��JПE�[5ɽ�*<e����@��F6�
���*�>�I�n���l�G���s�>���	2�B�'��hE���ɽ�*<e�ŕI�(^*��U���\Jԙ�% �f��S�Htz@L�A��V�)iɽ�*<eW�h;�A���M��ȶ���8�!�|ɽ�*<eW�h;�A�;�����Q���8�!�|ɽ�*<eW�h;�A��x�R�l���8�!�|ɽ�*<eW�h;�A��M�U�帶�x��]�ɽ�*<eɽ�*<e��U�kF�P=�ض�b�E��o��ɽ�*<eɽ�*<e+ֿ�n=��zȝ.�A	3AuF��ɽ�*<eP�7ٝGy�ɽ�*<e�+�r��y�f�{��t��
�9���򭸋78��@uk�Fg3�`xjZ�v��LMZ�"�9u��夣�P1޸��ϝ<��Uצt��y4��"���JПE�[5��}Gδ�-�HYd����ޛfe�^C�ɽ�*<e6pI�D��� d�^�K�m~�C��%q�q�����z�z�Z��v
�p\�Ì��:s��n(�a�K��J��	c�(��>} �J�rC�hbu:׈S�y��L��Ԝ�x���]L�E,4���?w|��\Q��:s��n(	���]��A�'2�O��d�^���4���?�ɽ�*<eB���0�|��K�`�r�d�X�m��K�`�{a�E̤�F+�m9Ku:׈S�y�է '������d��X��[��Ƹ�XS�<)�	!����M�|)C��:.� �0���%������ɥ!Tk�Y����~Q��ك�ā=d���[�M��Ҙ曥ח�P���C�/OA"��Yd�d)}�o4B!73G�,�x�u�o��'���VѐԜv�v\C�	���/��5��9�� ���j
6�#���؏)%�,�ɝ,����ň����S�l�G�N]Ե
Op�}�<[:� ̷�I�|��.��u�Wb�-�m, 4�r��K�7W|���!���F�W�����/�Q�t�:��ae�P��~�pԵ�l�j��Ǿ,GLY/E�Er�:�H����?�P*�փ��ɽ�*<eɽ�*<e6Q��f;��f2N'/ܕ7�D:u8�ھi��͗
ɽ�*<e��Ҝ�����%���x�aT��.�^t ��!�}ɽ�*<eL��*mZٝ�{M*�$L�pĹ�+ֿ�n]����zJ\bWM��>L�"۠��Ko��ԍ�E��5�l�dȚ]`u�D�ў�_bD����Oz�6|"��K����G���R�ʹXr�I,N��o+m��Fo�lS_O��k���,(n����67d���"���JПE�[5�p\�Ì��H
�owa��E��-�p\�Ì�:2ǑK��E��-�p\�Ì�Q��[1���E��-\Jԙ�% �f��S�H�E��-\Jԙ�% �>|
ϒ����E��o��ɽ�*<e+ֿ�n�Bkv^���NSad���H)��k��K�`��������8�!�|r�֏��9��W8 �+N��ߔG�=��*��ׅ����U������l�������&B��2���m�@|,�m�ɽ�*<et�%v�yWz���xE��W*X��!j�������M`.��>���	��\Jԙ�% �>|
ϒ���� �� ��Gɽ�*<e]L���z�W�D6�fg�IGL��(�I�.L;�x[���K&���j;�����p��O�
����8)�'�C��!DgW�Ǯd��``ط%|��r�Qx���]L�Eɽ�*<e��
����a�t2Ψmv�Bӝ`5��N�8Rlƫ��n),4���?wVm:��J]�~,��~�Ge.���U<1����c���1��gɽ�*<eɽ�*<e�H)��k��K�`��������D��aɽ�*<eɽ�*<e��l�G���/}�Ofgٕa��Spɽ�*<eT��%z�s����+��=0a�ꉂ�R=>pAJПE�[5ɽ�*<eɽ�*<e�my�odK��H��l��NSad��ɽ�*<e�p\�Ì�B�Xpf-��;9��S��A�Y��gɽ�*<ef�{��t�ɽ�*<e�Y�tѥEo�
�0�C�˳�Cd�2J��A��Ѻ� ao��k���,(nɽ�*<eW�h;�A�;�����Q���D��aɽ�*<e]�P�.�F��u�ǧ2��$���p2~ɽ�*<eT��%z�s����+S"C�J
��3/�})�޷����wx���]L�Eɽ�*<eo��Q񎑍�\=�6���Iy�ɽ�*<e���&B��~��\U�(�gƋ@�������p����8t�֨��S���?���'��%V3�-�Z�R�ؑ�JПE�[5ɽ�*<e�p\�Ì��H
�owa�dB��5��ɽ�*<e\Jԙ�% �f��S�H�G*�ag(DA�Y��gu:׈S�y��L��Ԝ�x���]L�Eɽ�*<e��
������������K�f��S�Htz@L�A�
���-9�$[|z�ɽ�*<e�_F��x�&ꬶ�R���&B��~��\U�(��5{�ѓ�͌r����ɽ�*<e�H)��ki��)~��NSad��ɽ�*<e�H)��k�F��ɱ8\�NSad��ɽ�*<e�H)��k?������*�NSad��'$��R��e�����kV�P�7ٝGy���8t��0.d�չ�RO7iB�wl��[��Ƹx���]L�E~4�R�T����/����U�������8��
l:4ʛ��M�x[���K&9*�b]���
/���5�x�JZ����qU��Oɽ�*<e� EOk��˳�Cd�2��/����`�z6ɽ�*<e����sMZgV�|��.LY��<0��������$�ɽ�*<eɽ�*<e�'�و����K�`��/�ΰo����7`�%���K�U���YJO���g�Hx��D��k�#�^G��ٱ�i�Z��?�9���ْ;0b5��u|R�2�i1���u�\��u�t���JX�o�'���tM#�/��t'���hX�O@g�IF)_d<�cYb�'����4�È}����Hc�;�Y^�U=���8��u������Qk4]��
�k���_=������Y�"�WZ9���u\�a݀P�!s�,�	���Π��U��~Hfu��Ԯ�΍T�:��S� k�7��`x\ `L����JmB6q~q�~�i7 :���Iy�;�nų�j �@V��"WP{Y�GT���8�Y��i����QQ*rbH�iA�UAKTnО�>����x�})I)���()�6��9w嚋.�����_xUʯfK���� �]Ե�:i��Ly�|y�ި���6�ʈ����I_�Ut�)��7�џ�q�s�Mv�'��X�)����qӬ�\ԗ������nx�I��	n���#���o�oi�8�,����̜�ߑk���g���>�0 ;��od<~R��Ǥ����e�9�\?%&�/�~=rN��uL�7d̈w�U���YEL8��L�Y���ay\�n ���J?|��'�[����K���3��h�A5�oD����S�_>gN0e�,F��Т�����[���ɛJ�z6Ǡ�&�ǅ���7�Y�}ފ	�c����$���D����,���AI'�Q�Oﴽ���������
����-��
�=��U&ʀeH��J�	�5!�`G$j`{�+!�Nh�z�{&�@�J˔Qm�4ߥ�B��e��G.I�TVzi C�"4D�ؘ����T7]���`r���"��Ip�ёg�L.M�"��P{�5�uk�]�ͻlU����\�IFw/�QL�L�e0�4��k19�"d��?0yB�ג$OJ�7��,v��Z����z%u=���a�ҡ����Sk�*;���>�v�E����>�d��xff�Z��>��(��dp��*��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8���ա8&�o�	rr��I�f�Ni�Q>���ě�T�t�g��g�����6T��;ڿwT���V���b=��K�X���hs������p��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eT#@�GNɽ�*<eɽ�*<eɽ�*<eɽ�*<e7��� h^������ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��q�Ӭg��K[%�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�S������k�L�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e���1Dȅ�J�_�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��!�2X����]��5ɽ�*<eɽ�*<eɽ�*<eɽ�*<e���&B��E����Ѳ�����p��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��l�G������p��ɽ�*<eɽ�*<eɽ�*<eɽ�*<ef�j�Kw� �p~rևD�io5CB�O���	�%�b���E�oGq-TN{��U~HɃ���.��k���-F��lB��k�9;�R]�������*���{�u���w�|�2a�3����o�����S�#��mIӛAЂ&�(�ă�R5�+ұ���_���G�C�L��-<��eh�V���tPfW�������)�orL�˝Ly5-I��a��+�~^<y���5��M���")p=_��ö)���')/�=i�S�>������yl2���� �h���΅�*�6U���-����S�[����~��Wɽ�*<eɽ�*<e��g]�?�#St�{j�6?���:�ɽ�*<e���&B�����|��.�Zr%����%5bڍ��q��� E���3T���O�. �������^�5�ɽ�*<eɽ�*<ecS�<�U��?��Խ�u
����.ɽ�*<eO@����,�JQD-���sx��f*��_��CEP�W`c��r���#5�*N�sӄ�]l�ת&��~�af��s�_�A��Y����m��c\N&��N��8�0����(�[�v���x}�IZ��V��:�N�c�;�X4�0͵�Fb���g�H3 @~4H�򰁓.��֖=���b@r���28��GB���K��G�>@V�S�~DYI�P�lz��J4�2�|ɽ�*<e��x�hd!p*�~�m���ZBV��9�p���h3��.
�_F��D��k��-O��V�n�&T ��c%�`V�f�Bɽ�*<e���M�����ӆ�澮/�žCɽ�*<e�^?��C�LS��i��8���'
���it�z���ɽ�*<e�^��"�6$xU�?��f*��_�Û��Uv�����p��T��%zؕ��g�q\��/�žCɽ�*<e�����F2]�J8�F2]�J8�F2]�J8�����p���VJUT���Cu*�Pf}��OD���Xyr5⊢`������{�:�0H�� �uɽ�*<e,4���?wX�1�{��F2]�J8�F2]�J8�	C7��3�^ɽ�*<e��}Gδ�-��~��]�xɽ�*<eɽ�*<e�?���q&Ȝ��X|�YA�Y��gɽ�*<e�5����fF2]�J8�F2]�J8�~�&T�S�ɽ�*<e,4���?wV�,��$�7��Cb _.T�!�ǥ���	���{����1͙�+my�ɽ�*<eZC��ʟc�r²�[���hɽ�*<e,4���?wX�1�{��F2]�J8�F2]�J8�	C7��3�^ɽ�*<e��}Gδ�-x�g�щȸ���������{|��S91��?��|ٯ��������ɽ�*<e�2g���VbD<_�Nɽ�*<eɽ�*<eN��-���"��FP�x\�����p��ɽ�*<eؼ��y^�ɽ�*<eɽ�*<e����jt�tz@L�A��V�)iɽ�*<e����,�4ɽ�*<e�+�r��y���8t������p����Yr5'4M���//�%
q�sڝ�o� }�uKO��m2T ��c%�`V�f�Bɽ�*<e���M�����ӆ�澮/�žCɽ�*<e>:�BLJe�����Ro��NSad��ɽ�*<e>^SH��⛱����Ro��NSad��u:׈S�y��L��Ԝ�x���]L�Eɽ�*<e�^ưVx}mr7��;=4Y�
�ugƧ)����ɽ�*<ei��y
�d,�
�a�ǆ	�U�5��/�žCɽ�*<e��}Gδ�-�M`.�ޛfe�^C�ɽ�*<eɽ�*<e��'�F�`!�׃>8�C
�V[�ɽ�*<eP�7ٝGy�ɽ�*<eu:׈S�y�~��MG� h7�!%ɽ�*<e,4���?w�7�T�N�o.XSG.�^b�Z�6�{ɽ�*<e��
����`�hP���^��/F.��ޛfe�^C�ɽ�*<eɽ�*<e+teM�i���^tD�����ߚ�V��X��Z������ɽ�*<e�v�-V/ߴ�aە E0H��r�dZɽ�*<eu:׈S�y|��5�L/%ɽ�*<e���)��<�y
��iV E��{Gɽ�*<eO�
����������w��#��+�C� j�Z��JПE�[5ɽ�*<eɽ�*<e���cXqM�3pI^C�����p��ɽ�*<e����,�4ɽ�*<eT��%z���@�&F��Q�m��Qɽ�*<e�ל
ϙ� ɽ�*<ec�֗�� \���
�ԓ���i��Yr5ɽ�*<ed ߥdw�#w���ÿ1l�XiI�����p��ɽ�*<e�Gx��y�� X/W�6�61MZ�SY�żɽ�*<eɽ�*<ei`�iWӤ� j�Z��JПE�[5ɽ�*<eɽ�*<e�ݶ�<C��M�3pI^C�����p��ɽ�*<e����,�4ɽ�*<eT��%z�����[K��PM���iwG�]v�Q~gƧ)������8t������p�����Ɔ��"H<��T�wp���	���*⬒��.$�K��G�>@V�S�~DYI�?��f��h~�L{�3�"j2�����+2�`�C�j�o��F�k?� ��D�A^?��M��z��R���{{gy2#�
R��r�=b)?��t^��4c��	ko���5���?^� .	��6���TXޔ7�ߞ�9|�GȆ�v�V�W�v#@CH5x�`{ѕ5��l)Ȟ 胨Rʮ����=����M�����ӆ��z�wjr����jt�����չ�<��̣q>Β�,�P�DV}�N��#����wW������n��4R�1��}Gδ�-�F�W����ޛfe�^C����!�@W�s�>�����)m0�-�P��^��x[���K&;������W����wW��ݶ|�N��J��LtE�����,�4����0bH�sm^=E��Rx�r������spoz�X�}��R��Z�J���F�c�q9r�T�?:�;���A��#�P:\����u)�QX^�2���@i"M6f��������5��	"	���?��o��N�1�a�g��ۓyP������1��
O?�p٫j��"�yL�x���Ys�}�q��?Xٵ��5�,����F]�J�������	UQQ*rb�5��6��uF�p�	_�P塙@:/!M_[V�I'�
n� 70^�d�e»�-0^��,�:�	S�uP�M�zK!�g٪�'�)��F�p�	_ى�#�9�$�oWU� ����L�m�C��#��;����B�	?�gwC�N�O�lK���K)��F��P������_#Ǚ��R�����'c.�	?0-� ����Jv���,����@p~�@oH��{T��qɮ����D���,%GJ�=�rW�K�v��|�5������zWG����ʙD�0@]�����>'�6�*�q�t������ϩU�R�4�t������:Wp<!���I��d�>�r=D�9�)�Ί#|�Ӏm��!Q	s>R=��@�wG�ɽ�&���[�O�VG/"���@V��"W���à\j����f���ԝh<K��}|�?�M��\%i�������E�!��o�8���RX<���O��"P)�6�m�`�� P����Y6Z����*y����,��/�&�5K}�*���ՙ��e'�������s�SŠ��z��Qd_No���?�%6=��� ���z�ȯ����2���Ե+ĳ�)[�AM]�찴�}0����:6g�����6T��;ڿw�p -����b��i1��i�y����4\��]�찴�}0��"�ԏ
�}#8�mÉb=��K�X��u�Md�;y<�ZX���}Ո�,�AQ]�h�j�v���� ��B迅9DԄ�r7uo)V�&�>\���^��0*e
�Xne��ƍ�C��y�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S� h�����\��^�9�>���W�n��)�p��3Ԅ�"��Ip�ёg�L.M�"��P{�5�uk�]�ͻlU�� <�ZBg\�u�<T_?�O����X�_�W�_�U���Ɔ[����b�A
t�Ke�%zQ�C�L��-<��eh�V��KdiF+N��l V{���Qv��J�Hw^���r���Oi��%~���m?\���cWΰxQ��ƛ��W b;~�1�ol0�5�s$0�D�R��z����%C�P�>{9pI&(V&L^����d:�yPl5uK��!�a�kea������yB=�u�@3��g}Z���O`���}�{H�������̱�Hv@�����JY�?�4h��p����	�:����8!��ɭK��7~ϓ��;�&��y�2�I����fR����̚�RJlJ��L/�>b=��
��Z�8Q$�+���������%�5�;u,��7~ϓ��;�)��kT���~FǙeB^��r]�Ҽ�w	�x�Ae�+Sٞ8���k�ֲjx����Q��5��Oh`m�&��l�G���R������HY3%H��'P'���J�X���	玡&��!Q]�VF�N4��>R}9���7���ٗ������|>��N����"����mJ���M*��K�`�"����ٓ� l9L�8s6��Z�hL��sk��H/���q�X0�Y�P��y�C3-j4�"������_���G5�td'P�TT�I��~��W���q�ޤ7U*���g5��Oh`�w6�-���u���e�yp$�g>���|>��N����"����mJ���M*���3���]�Ҽ�w	�Y��Q�kE�ML����W<:K�#����G���R��h�!��qӄ�]l�תiZ�zt)�#>�����yN�F�8I���W<:K<��d����͸8yw�T�>Oʏ]�i7|2d>7'̨�p�k�r��s��
N��p޴A�h���f���W<:K�n����\����0TC,BP�/��u�g**��]���ѡ��E���I�e�$�g��t�ic��ݤ���V�+G5�td'P�TT�I���W<:Ke&����h�V8��+ Z؋$��,!W��
{�m�Ť�ɡp!�����E-a�͢'̨�p�k�r��s��
uZ�i��9{��������ow����2Q�-��EQ���ߕ7~ϓ��;��T�vo��%H��'Pt2�S�f��
��Z�8QZ ��R���s��~�L�����A�>�����z�_���F�y����4,���#�
���F"x,��/kr���2���C�sNq�0a��<	mꧢ��O��xx�_x�'��4�2��R��얰�s����|>��N��a!�R �\�H
�&�0�@��'>�ԊȜ��X|�Y�֝�%��\F9�l�G���R
eka%��A�
����eU�h�-� ��׼5��hm�헃P�� ����y(���f*��_�E�I����	td���AgWf쎄X��X��ZC��)p8B���7��lEX�A�.D�K,�%��5���K��������� ���������x�h�2��B��:��� j��!��ɭK����é��U�
��'����<	mꧢ)� �)X�h�[�E��%�[�R/��w�#ۨ�D�_�̸B���3�\��b����<���^�0)�D��+�r��y�z&ŎlN�/��t������_�%˝�=��C��e����>J͸8yw�T�ޛfe�^C�(��Î�HX��	ko��-�U��8����p��mIӛAЂ������CK����=��ti+L�h�,�B�iZ�zt)��Yr56����S�WJX����0\���w?�[^�l~%��K�`��_0(����i��g���V׉�1I�8[��)_�\#���aI�����DE-a�͢�q��G8�i*3ZC�q�����w� ���x]��ג6����S�WJX����0\��u�2��] yB=�u�@3Z-g4.��E-a�͢'�������p��mIӛAЂ������CK����=��ti+L�h�,�B���6��F�G�8ٲ�X?c6)ܰnslf�{��t�_�����l:�!�@�5�{���rt�˝�=��C˯�C`�*֗�s9�鳓JПE�[5��^/a��헃P�� ��xȭА��f5���c%H��'PS>�tv�x�O������|>���qa͸8yw�T�"䀊��Z ��R�
���F"x�<	mꧢ)� �)X�h�[�E��Z ��R��e����é��U�>R}9����é��U�����z�w?�[^�l~%���!C�P�7ٝGy�����/ַƭ7X>�їT�t�g��g�����6T��;ڿwT���V���b=��K�X}(�K�r��ԉ�O�F�ud�^jN�z/32]|��JR��v6�![������IpK!�R�Ժ�:������M!>ܼn�xQ��ƛ�խ:���xQ��ƛ�0Ȉ����P��!L�c�`�eg�g-9�a��M��M!>ܼn� i���C(��3WWC����#�Nb��PAv�'�B�n�Q�]��/\2�<MW<�M`.��M!>ܼn�Aiq��%���I(����A����#�����\ցKB��"3�^�&�������*>|
ϒ���+�>���4��d�B�:Y���!����(da��E�� ��׻���0�(��ݴ��D��{�w�Aj@��g��,i0�X�)p8B����9��V�c7��g�+M�(�bJR��S���� ��׼5��hm,�a��@"]˪�ߖ��q)
�/w�Q��ۿ<	mꧢ~�����Xƻ�2��x8�U=�z���V׉�6s��}��L�<y���$��D���Z2����/P�c��x���]L�E�(�[�v��>S2{���G5�td'����4��V��P ���^�W�n���Yr5���������y(���f*��_�V$eHIĉrmF�A�*k܂0 �f*��_��{Vent�L�"۠��JПE�[54��!��	���jq�4)0���L�m���f���n]{�/P�(��Î�HX����V��ym��A��F���e&����h�V8��+ Z��1�L_��_0(I4������z�ɯ�6$����>7�(�����\Nh;wݧ��n��� ��몊|s�=F�`V�f�B�j�8]��{�w�Aj,�o��v���0����xȭА��f5���c%H��'PS>�tv�x�O������|>���qa͸8yw�T��y�f��ɽ�*<eӄ�]l�תlL=L<[�'���D�cQt4dB���{Vent�L�"۠��JПE�[54��!��	���jq�4)0���L�m���f���n]{�/P�(��Î�HX�m��c\N��K�`�A��K���ɖY׎�YZ͆ˎ�8�K���V�f�o0�$���<b2߯AaI�����DE-a�͢�q��G8�i*3ZC�q��`��$N�+�����&���0����xȭА��f5���c%H��'PS>�tv�x�O������|>���qa͸8yw�T�"䀊����|>��Nn��i;C}�Z��Ct���f*��_�V$eHIĉrmF��:�1Qb�ꔻ�K���P��;���ɖY׎�}�tؤ�l�k���,(nWCN�;������%�;��\ÑN�wg�	��%���@����^/aË(t��S8|�t*lC6t���y�P�+�r��y�z&ŎlN�&�	��o���?��h;wݧ��nBP�/���/P�c��x���]L�E�(�[�v����}nW"Q�����4d>��q)
��:��� j��!��ɭK����é��U�
��'����JW�0���~�L�����3�9K��Ť�ɡp�:!����P��H/���y�f��ɽ�*<eӄ�]l�תlL=L<[�'���D�c���NZ$i7|2d>7eV3���MJzA,��geOP��;���ɖY׎�}�tؤ�l�k���,(nWCN�;������%�;��\ÑN�wg�	��%���@����^/aË(t��Sr�qr��/_t���y�P��?��zF�	D�ܣ{U�荑Z��3������Uj٨ꩍ��n��yO]�&��I���R��A|`�$������kȡ�B,ŭ_
j�����ͬT$OeMS���s�C�罤�9.�f�i����
D��H7����{�ƥUuh��V�g5D�l��9q�X�:׮�5:��KL����z�>�4[���{u�^ק��}�{�ʘ��SD!��Ю���0�V�٦�����2���X�����wD`֡��y����"�m���F^��`���#H����^'�2����:W�0s�����S�_>gN�-�:'��$+���G(����^Le�0�[��z����jcbb_�B�,��y8f���B6Km���'�5uEq_�<|7.���|N;X�^�I�[\o|�o�����|"ÝW}�utiO����+�%�Q)=d���E,��h��DZ�x���F\��w�0��8w���c�Y�l�%�tB�*��� �&&s�:v3�9?k����Q������L�����p�N_�qe�
��>̊��%�
�T���k���g���*�F/��q+�\��$|?G��a�G�x�D�9ϑm�eQ���9*Q����� P�7+��$-���G[�z�A��ie�\#�_Hc����'d����uC)�E���Q�0)Dm*
kma��ݑ�`��N��X5/�)I�|��o9�H[��UF�n]h�^�o��p����=����+P
���(�5;B�W��M��v��E�`�w$�P��j�:�mheˣ��:��?Dg,2ms����{Ue#T�U��nl�ɀ�\�����;�������G��Q����9��
-dϦ�}��0�`�+�\Z6��v6|�d"81�r#���dxxoM�L4ğrF�}�����'7�{Y�R]u�F�p[�:N�Ƕ����{*�㮝�O����8-��AћZlϙ���7��AvO�:��}n���d���a�|��H}T=!�1�((J\$��$���Z�^?4�9l	�s=���fG$�8�#c�X�����r�lI-�-�����q�����[�p�h�-��\���8���B^����`�Rzt}a�Р�m��X�]YLچ��6�oє�B�qkq��x�`�K�[�!�4�9Qrc�*��������c�����t���ݬ��0�`�+Y{G�T|r>�,�L�N�#fH����2�&�o����6�xФ6��4tɛY�(��Q �:���2-|g�����l�����2-|g���W���p��W���p����  Q�#�|�O�3&���uL����K� ���ɽ�*<e>X����5��"N06F����/�N���JP�����L7bZem�ۜ��
��i��ȿ0�����w����5����k��$È,������Z\��s����Xg#~yj�FD+?��E#�����'7�������vTX���}0���6uĘ)HL���+�������7R�1��l�\�_�	(��X*?�A��jx�I0獰H�tHF��#��g:�Bح������A	s���B�p��3Ԅנ���Սy�ex�e��j.�qN8~N3�b��i���sX!�t7�e��cAe����]V&a;Bp_��r�wЄb��~'yE�"��Ή�Hh�t?kE�O�"�tZ����]6�[8Iol|e��j.�q���I`s.���$�P �Z��+�yoCD����(��e����� ��#*&h
�<�I��¹�� ��'f����� ��#*�E ���X���?),��5��M����h�M̻��wЄb����)n���M,�Q�.#����u��
�W�+�g�����]u�n�L�ߨ���H�Z��c�x4�(��r�����v��w��Kh�&�B��e�̣G�vSo��¹�� �=Д���v	!�k�$R�
?�	��%V��ox$���\فN�ʆQ'Ь�.e��V_���#����}�n���/(:FՓ�	�&�ԃ_��
?�	��9��1���'B��E��;���l���#��ǎ�U�#�.����p����*H�x���V�uCM���˺�1V[�wNʷY�rE�[#�����:��P���wЄb��':�8a�S+�n�/�GDQi���0ʇ��t�i�9�%�����P���/J��H�ABL�\��-���蟣��B�3/�.��+�>���1AiD��D���g'ë���{�?����޺��1�0.�h�+�C�.�B&�M�3pI^C�Һ��F�YgƧ)������.e��V_���#���;UT���2�[�_B�|'��v����aY��ST �Ǽ��ܗszЕ&��|JПE�[5C7],ρ��E����k���l��H��/p3���X�aҥ��)o0$g�`a=o���
(-��
�)�܌>��<��+ʇ��t�i�9�%����'f��ؼ��y^�p��ۥ��}6�[8Iol|e��j.�q��a�D��(-��
�)�܌>��K����Ɇ��q&�:��R��ȈGn=�-���y���S�ӗ=E��Rxx*ّ�9 �#P�o�E� :N�`�+1�;ی��gt����%ZRh�U�*��nm�E|�N�)��A�Pɔ=Y3+׵`:y�Z��������|�����N���Q�)y�˕N�*��3M>3���2+k���.��W��[ݬ7�_�� ���	/�2+k���yN�F�8ItGD���R���K��W�\�.��~]��K��W� ���	/�R4�&%q�*9�����DF��t�1	T=��q�77NO�����DF��t���q�>���� ��:��;����dk|������_�ޔ�~M�
�� ���%6�G޶���-p�!�6��q1���a->�d�wo�	h�[�p\�Ì��F���T���a->�d�wo�	h�[�p\�Ì�46��v�k~ƅ=ht1\�I;���ɽ�*<e�2+k���+�(�T	���~��WO�"��Ǌ�7�3x���O ��sye��yl2���ɽ�*<e�K,V[dn�QD���~��Wɽ�*<e�����`��\�.��~] ����E�.�^<�
:�ɽ�*<e��X�Y6�s-\a�"G���x��H�iˠj&!��E𭨶H$�W<(u
����.ɽ�*<e}!�Lڜ(,�QhfB��4ud��E��*��c����p��;�Y��##7�1
����e�̣ɽ�*<e�K,V[dX P��>d}�v����O�"��Ǌ�1�C��~��1�A)��2Sn섮�}>N��W��j����t.��d����H<l �K��G�>@VQ:%~$�>%��}�F/�zo��&�{NcB����'��`
z�A��(4�3Gbl��� �&�-1�>l��[�^4%akԅ����	�\�Ys7��Q�:��})~&�X*�wЄb��"��:s�8�uh6u�<�]�ͻlU�� <�ZBgy����Q�%D�M�Vw�ԔD����y��Z�ՠ��sCܛJf,ٵ����g�v�\�`TCܕ��cWκ�;?Q3�q���o�(]�}g��+�n�/�G&h
�<�I��¹�� ��k���Z�8}�Rk��k,�����p��l����x���BFh߿mh��EP$�"Rݗ]T����R������֍`,-�jл��ukԅ���:)Ɣէ��Xr�߂���q�E�Sga��&M����Do�3�uѨ�<��8P��c�C������o��������rZ��
YL����4gT�d����L������p��=F9��V�TO��B>(�k�$�t���y�P!ՠ��s��Y����Sk�k�9ע��Z�k���8t��}�tؤ�l�k���,(nf3���W��Z�8}�Rk�Sk�k�9�Lԏ���6;��2��:7����@��a�N�~%9�t<ŕV�(�x���]L�Eɽ�*<e�n �u�HY3�P�^��,{sm���8�d�	��ɽ�*<e1��0�n
�(,b`e2���n
�(,%y?�>J�T�ٝ߄��s8���F���'b�$d?�Wޔ-�R��-�|�L��y�wa/1�J�[+S_O��k���,(n-��ó�ڋh������>���o��3|Q}�{$��~-y7{E�6��h#���T��/�����7R�lhL�ɳ}���A�Y��g��<��ݭ�`V�f�B[�Q�X"��|��_�ޔ�~M�>���5ׄ<�WV
v�,��O�	�u����Ɇ��q&�:Y���~K��ٴ7����~��Kn��|�;�&�Ѻ mT�AMu:׈S�y�է '���x��D��k�h����5\�YuW��<a�SQ�7�Xd`�,n���!���8B`}�'�4���[\�u�<T_��֍&b���gc#��ό4j9�>�u����3�!X�Շ���Q�t�fɗK��Loح\x��?B��O*�*�����p��ɽ�*<eɽ�*<ex�\�u��9��E�e�$���;�
g��^\���q����5L�M,�Q�.#����h�	��_Y�o���n<��4Hw^���]������˧YR;	{�_Y�o���n<��4Hw^���]������˰U��A�>R}9�ܕ7~ϓ��;�u6��(F���=���i����Ȟ�Vw��xZ����*�r)W���9�yl2����ar��Z�.�_7"<Zr��"�����sʶ��6L&ꬶ�Rȃ���p�����N�������Z!UB+����5��Oh`B�VT�́���b�6�}<�T��z��� ��#*����Z����m��h6m���q�_n?�?}��~��WRKD�vQF'�BI��^{g����M���K��-x�yl2����ar��Z�.��n���=�W�^a�ȧ���/]�Ҽ�w	�I�D�J�:j���+�Xq��hH� �ϵ%[��zN�����R��z��#	w�0u�a� z_.?�P��Y��G�y	J�X쟋�yN�F�8I���W<:KRKD�vQF'���_<+��c��"�����sʶ��6LycxB}��ɤn �u�HY�(`h���w�)3��Z�������NX�Jj�*���k�L�����N�������Z�2+k�ݎ�]��5�5��M�����x��{��_��l�ֹ�TC�r�r�Zjsp z_.?�PZ�������%�H8�`��N&�=�����W<:KRKD�vQF�z�H�?��� ���	/ic��ݤ���S���)�!ɉΔ�D@~�L���7�'`� �����u�i7|2d>7��M���9-��ǿ�B)b> |�!Nic��ݤ���S���)� �)\I�[{���J�n0��?�Π���Z��G�M����(���_��{n��/��*��0϶���;6U�l� >��u�<�W�~��T+�ͦ��"`1�t�~���O��m\Ʒsa
�B��#�c>�����8�À�؛w�4���u�C��䕊�R�NBQ~[��*c��ȥ������%��`��-c����+z�%zu�Z��W�պV��v�'�8wnr�����r�w�|ћ���|s{k�����)Oa��zu�,m^$cI�yڡ���R=H�q�b�R�f/�V��n6?l������:"��
� 쎤d�w�r&+��1dQ�On�s���99���n9Ð������[(O������E����R#l�>h�t~&@m�`+�?�nr�������D�����Z�D��������)O@��F�ZO-1�>l��Z�����ų�J�ٌ��T2�מ4#vJ	M��S��^�
&��bM�^��_��K D6I���ɥ�ZKϘ���F,?G�i�G��}x���Q�O�. ���RKD�vQFEŝ�h8}x���Q��+�(�T	㠎{v���su�GA���O<�O2|��ö�#5����Z�O�g8L}!�Lڜc-��Ο��zN�����66/�@�H�I>/�4	oZ���E��uc�逭�p�(�4���Q'�@��.*l ��55v'��m�O5zws��$<Q'��Y�y�����2G��V���L(���5��lP�3h�4����uhN�V�Y$������֦��u�j�+:4ߥ�O�"|	���VHU鄇y��k�C	x;�����!��d��M��AJ����§���H56�	OƗc�p;h��rRo��b�;lly��;��`�A�p96� I���e�ιv�����1b�_or��QM�f]9�A�H��;�s�55v'���r������>�N�?H'1LC6�^��_�Ϲ�%��09�*��(���FC�1|�^��_�ϕ5���>�a�X�%9�*��(�b���ƄcDr���M��ح7{���V�(��$h#h�¥�P��`�a�5,�-8�Y�&�9\�&j9D�m��I4���Z�۬���-�.�t���%D�M�V�5�<z\u
?�	���3�T�JS=8��d}���p~	B�+�n�/�G	�y��pW���1AiD���cWΐ>�g��kd�WG
�� f�Æ�=�6\%i���7d�"y+�7��Y�5��y�)�\y��(�d�� $��f�Yv���wE]�ͻlU�� <�ZBg+�n�/�GA! �+Є��?@�����cW���cE,j�0)I�P�z\�]&/���_Y�o婛�F��K�G���cW��p&��/��Щ.�v������p��ڭ�b�o1�`oXO&�Jڋ{/TV�x��}r!b&X͸8yw�TيUW����yB=�u�@3-��F��٤�`������u(t���
��2ˀF���x��ɽ�*<e��D{�I���V�uCM�����jɽ�*<e��$w�[���V�uCM�b���o��ɽ�*<e��%Ho��^���V�uCM|�9ryɽ�*<e�T�g�lsq'	�7�G�'��:eA�9�W�^aǯl�SX���S#��\���V��o���V�uCM������h6m���J��E�i?�W�^a�`Z#�V>�����p��- Z��(����l`.��/n�����h6m���s�qRC��:+�n�/�G	�y��pW��<�{C��NYD1F��Y�rE�`��%-�E������{6��SD+�?M�Ȧk�v���v��̟�}+��c��{6����hƁ�,3D>�d���q;��3�~7�p�<$��儙'1vdf�f�+�n�/�G}!�LڜV�wX[�<}!�Lڜ3D>�d���q;��3R�%�v�s����hy�O͗�^7_�ŕ��cW�� py�;�PlS�������k'�{+�n�/�G�e�4Z�[vQ1��􎖃�1AiD���cW��V���0����F�Y���A���t&YjԷ��Gy6+�$��B�Ơ�t
	��f��R�P�y�XX+�n�/�GMh��A�Yi���zT*�a���+�n�/�G)��¹u)^R�m�J��M�U�帶J����A� L՚`Rp���yɼ���%N,��t{e賙m8E�G��_|ѯ
?�	��Q��	*,#�5	��j�S�ح7{��'H==s2��_o1�1\�$���P�8k���d�VO���]���,G���B�S�K
�
'P�4�p����4\��]�찴�}0I�cl�����=��(P��q f�&�����������p���'-�rEJ�H���vN���+����wcU �(��K!�R�Ժ�P��a�'���cW�gSr\B�Ԉ�*B�qRB��2�ȡ����$'3Z�R�Ρm~��c/���Y�G+�n�/�G)�o{6f>xS�u�c�z�#��gP���|s{k�����)O�#-�g�sʼ�WJoLg�l'N~�*j9D�m�����w�x;�v���9� =s���G����1(a�q<��[E���V�uCM9�R����q(0)�J��DS&63�� =s���Gy�Pd�T��z�`u�t��s禩���`���2�ڞ�up�� b�����V�uCM�UopfU���	_�������p��U�1����Y�J�`�9��H�Br��f	������p���<�����=+g@{���;�Y��##���V�uCM�#�����^F�4���f,E(�3r��?��Up"C�U �>|
ϒ��ޣ�/��O�%� b�������m�/(:FՓ�	W��<a�S�R_t���P�O$*�ג$OJ�7�-h�+��y����Q�%D�M�V�{۪��w��&Cx�,��'���*�[T��/���w4���xWz�j�+����p��!��l�G�p~	B�+�n�/�G�;���J�z/��[�Ţ��?b���1AiD���cW΋*,m����Qb˪0�V�u���ᦲc�����p�������X��VO��۫E%��D�&8���í�2"������Ҁ��y�و5���@ԀoT�hl؎�	�y��pW���1AiD���cWζ�>B(`:�@	 ��U�+��c����V�uCM��c-������)|�RW=CՂ�z���o[�u}Rk!��<�lZ���,��(:��	�//:����#�>��xl�(T�飳������?ʌ�of�F��i��e��}R�|��W��A��1�����k{��Ty}�zj�"��0��U��j )���.s���2D��%_�y��N�[\��NT��>n.r�P�S��И]h����,��D�se��L���Ӡ��B:l��9q؟��?��6\F�߉�}3z�s"P�A/5���{�)J�ɷ�b���Ւ�tU#�݅�Cs����myW2��KqM�qsdu��&� �r��j%g�*E�Z��(wRET�1�ZAů� ��Ö|�o�l&��H�J�9B�ˎ�U�X���!4��x�ٷ�?��Ŵt� ��R����a��'��FL�j�4F�tˎ3I��(��Hk�p�IwЈ�#oԓ`��Z���GD����4�fgHg)%�RPz
2����$_�>U�V�Q���L�˷P�B�p1����Z��U�`6�!R�4�t���!���8��`�w$�P��j�:�cb�S���mheˣ��|>X,1��>�5T�g�'y{�I��y3AL�����~ָ���}R�|��`iX��-�����I���#^2�}G+�����uP�M�z�ڽS7��v�����
����%�z�M	!��Ɋn�]#�$u�	8'x��)�)�����y�>�t�Jд��߿Kv���������0���L��J���n�+cb�p�f8��H�\=҉7�#�?hX� ]����f�y���Wt򐹸���9l/-��փ�[��ў��4�IM� ���	rr���6�XoND�Zh��=')��ˎyN��d3M6�J��Vɖ�5�}�'ҡ���TX�G��Sb=��K�X���hs��x��v}e	�qu8U����t�e��*�Է�Ө�wO���ˎ��/� Q_�ؾ��S#��\���V��o9UX'yI�E�TҘ��S݊&�S_V*Nq�t��|�W�^a�J��^��@*Nq�t��|�W�^a���1dj��*Nq�t��|�W�^a�����-�'�BI��^{g����M���K��-x����m��h6m���J2�֌�!���w�2�(���-��@�)�R#l����S3.
ꢕ8�'��x�=|k�^��r�rz��� >��	��
�E�&�7Iy�.g���'u��j�+N���+ ��������XVt�m"[°_�w���ʌ���߯,��"�e�$�s�XCjf���7��pÜ6�w:�|����9�ִ�u��_����R�bT~����<�����ġ� ���_Ʊ����7#poGS���д���W�X'�/�=,3�2�(���ܴ|Y�f���t����{g����M����%�{W��:j5��TҘ��S�n�T�g*Ֆ �~o�	[��ݒ�J�N�jw6���]#���t����{g����Mhh<�i;�{W��:j5��TҘ��S
r���t��?�;D�m�n;��w�h�r7��qz�rیm/�=,3�2�(�����V�3�~޴	�E2}���bf�\c�=����cq9�toDTS�����/B	��L�fG]���eJ�y�T�������D�~�;5��q���T-^�R{�x����k�.�����2I��	W\�Y�r�O˖1#���p�Exk������2I��G	��F���w���y7�(��#��$f�A�$8�Y��L=W�x�G �����E��r�pRZ�r��jf��@�'�^Y�jG��Y����W�à�{v�����X�?�t�Og�V��@:RR�5=�Q�w_��T"�9u����'>�^�uھi��͗
�3Iw�cG�LL�1������h3��җ�?%��[[$6��B��Ę�c�����:RR�5=�%�4�5�V�\~_���c̘��V�!8�IF�V�\~_���c̘��B���_5M[�ʛڪYɽ�*<e,�x���m^{�4r�~WƱм#�ɽ�*<e(���X�Z�#�Y��%����cW�ɽ�*<e)�I�����'>�^�u���V�uCMɽ�*<e�����{�
��v2� ɽ�*<e+�n�/�G�h���K:RR�5=�G���L�w�ɽ�*<e��:eA�9�W�^a�	���!�Y�n;��w#7JK���ՠ�q�1�ɽ�*<e��:eA�9�W�^aǓ��"XH�nn;��w,�}NhG}�ՠ�q�1�ɽ�*<e��:eA�9�W�^aǜ���[i�n;��w��u7<	�}ՠ�q�1�ɽ�*<e��:eA�9�W�^a�Y{0�h�;�n;��w� �g�e�ՠ�q�1�ɽ�*<e��:eA�9�W�^aǤ��q�B�4n;��w ����7Uՠ�q�1�ɽ�*<e��:eA�9�W�^aǨk��Tzn;��w�h�r7��ՠ�q�1�ɽ�*<e��:eA�9�W�^a���B�|���c���M�J�N�jw6�,�� ��ɽ�*<eW���P���S#��\���m�?��i�����Uh6m�����d���>ɽ�*<e�VJUT���wۛփ��A���ƍ�sv�{d������p��ɽ�*<e�r�`�7ɽ�*<e���D{ V�xf���cWSE3�	čɽ�*<e+�n�/�G6�O�C�8	���!�Y����V�uCMɽ�*<e���D{ V��J�N�jw6�)\���Y�ɽ�*<eɽ�*<e>�Z�('����D�0����g�N�kɽ�*<e�����©?� jLⓊCU��eq�����cW�ɽ�*<eq�AsףMX:��/�M����Q�,ozɽ�*<e+�n�/�G6�O�C�8���"XH�n���V�uCMɽ�*<e���D{ V��q͜R*��Q�,ozɽ�*<e+�n�/�G6�O�C�8���O`ƃ��V�uCMɽ�*<e���D{ VΨba�dQW�SE3�	čɽ�*<e+�n�/�G6�O�C�8��E���W\�5oҳ�ɽ�*<e���@�-	b=�(|�4A���D�V�ɽ�*<eɽ�*<e>�Z�('߭[M��hp��g�N�kɽ�*<e�����©?� jLⓊC�&�K�'~����p��ɽ�*<eK�T�L���VV�*H���g�N�kɽ�*<e�����©?� jLⓊCl����&����p��ɽ�*<e��#�~I����p��ɽ�*<e�ޢ��X�[t�Lq��O��]�Q������ɽ�*<e�Xr�߾|�h8׬\"����?c�$��!,�ٮlP~^?0�����[/���7#MGʹU\��yJF��A�p\�Ì�V�\~_���c̘��B���_5b��RI���krC���i�eá� �)�[�Nz���d�O�,�����\X�HDč��D��A%�w���?��������p��0c"�&���N�Q������ �Ur��rQ���EP{3So_����T���,@�'��,���˨[�Nz���d�O�,�����\X�HDč��D`X�����7%�Jsc�RK�HxW��ʺɽ�*<e��3��c���8��i� |�oR��kc��O�V�EQ,+n�	��[���-����u��P|Ý� "�K����KE�׈�P������$�R�"SBe�;�ɬy�H��
���Ý� "�K����KE�׈�P������$�X�H	>��&�aC�5����cW�c�$��!,�ٮlP~^?0�����[/���7~�(jN���1�j�8�x%���%���&ZtP�S+Do�|dd'�)��"��Z�ٴ#�����4i��7�4��V�t4��x\��斳�-S?l��;?7d��4u9{0��%�Zݪ+iLr�hNev5���&���H p~�(���V�����;���03tή\�t1\nr�����Q�}c3�� �ߕ�"�;xc&z�j��S�#���:���R��K?���^��=c@�LT�]��rF���NÃ�u�D�>Nn��?_C��jtɽ�*<e��UMK��o�8�$7�B�q&os�'�)��חM���"!RW��ODA�Y��g��x	���8�$7�B�q&os�'�)��חM���"!��5;ԭJ�{�;���Ę�gu�n2�6�}����uH�������Y!�aa{�;���Ę�gu�n2�6g�}�zLW��S#��\���V��o��`?�u���^/a�61�fS�7h6m����
No�	�p���p�g�}�zLW��S#��\�ll�����"��"F����?5ǳ:ә�UK�W�^aǑ��a��4i�"��F�+n`�4"~��<ҝ�+�H�&��g��#E�x��*��~������#.?��z{�;���Ę-5��۬ɽ�*<eB��,Gv-;#^s�<����p���<��J��Uȡj_;p\"��K��f�{��t���:����F}ԥ�+w�ק��J��;�)>-�<�A�Y��gJПE�[56xOHx�R(�/��"6ӄ��PZVC��V�+5�~��`Dt�A�Y��g1��0��%���G��.s�x�c�^V�w����:�x*�w�Z��p��޶(:�`V�f�B����@��y�K��8�%aNe߯�-����p���<��J��}�o�$���8t���ɖY׎���ULf���DY �5�B���è��쐾�x|~�]��[��&�������p�����5�M�JĦv��ɽ�*<eg4�g/�W�릣� ��P�7ٝGy����J�Ij�2׉��N��gc�6p�h��<2L�?P�t����޶(:�`V�f�B����@���oŘA�Y�OAkHyaB(��[�YB�:
�1?�F������ś+�r��y���� �A�s�m��!�H�n��[���&$9��P��h�����޶(:�`V�f�B����@���H�����͈�3���ɽ�*<eg4�g/�W�릣� ��P�7ٝGy����J�Ij�2׉��N��gc�6p�h��<2�e*U���޶(:�`V�f�B����@���Z�����M���B��B(��[�YB�:
�1?�F������ś+�r��y���� �A�s�m��!�H�n��[��(�3�VE��H��*7 ��!Jx���]L�E��u�d�J�Z�T��3�*�6}�'}������fnj�K�P��mW���I:��A��K������p��/�%
q�sڟ��_V�c��&Nꊓ�H��d�
���WKRə��.U�[�x���?� ��8b�I����g��#E�x��*��~��������Bv��c�'�:�����W�#Ɖ�A4>}�(�o�%9�iK��A�Y��g��>O0���\!����JAiQW����P1޸����l�MojP�7ٝGy����J�Ij����W(���c�^V�w���C�
�l���^�{�
���|H�Pk���,(nQS��Df����׃/�=�k�)�bW�=""���J�G�`��ƽ.>rm�-^�*���|u��^5)��ɽ�*<e�V�W�v#@���M��L�u:׈S�yB,���m��H,,���c�+n`�4"~L��>�t�O�o8��5�1��厐��&�������p��BP�K��Rb�[]5�oZ��%�����o�����z Rs����p��4��z�#�t���y�Pg�k.X%1���<+Q_��|����kf�{��t���:����F}ԥ�+w��<��J��}�o�$�V,L��s�Ծ�/�žC���)�
4b�v�60�>v��!�l�ۆ�N������G���d��8t���ɖY׎���ULf���DY �G��<4b�v�60�>v��V,L��s�Ծ�/�žC�`j��V_3�*�6}�'}����4֊0�� 2U)e�YJ����,�4��;*��P���EXP(��e7�Rj1@��pO��'�8���F��7 Z�ˋF~:t�A���0{����&B�����9���x\gt���:u�M�*V,L��s�Ծ�/�žC�`j��V_3�*�6}�'}���� ʅz�)M�U)e�YJ�*���|u���x}H���������!�l�ۆ�N������G���d�CVE�OjN8��%q+�/EI`h��	�Z�S�s�+�r��y���� �A�s�m��!�����k�Y���$�C����8�O��F��7 Z�~��%0z�����b��������]�P�.�F�f�[>��������,�"��c���#H�N�}P��JJ��1�Ժ]'E���iW�C{j����kF;�x��*��~�������Ɇh����˖��.?�pS�rX���ɽ�*<eJПE�[5ɽ�*<e�=�ƈ���3�e4y��zɽ�*<e�r�\�׵�\N>�b���/����T�����1�W�C{j��뤫iga�Y�ɽ�*<e��^`�/�s��|�����lHkd�&*�]u��A�Y��g����,�4P�7ٝGy����J�Ij2�b�M���[n�+�'=E��Rx�+=�&���spoz�X�}��R��Z�J���F�c�q9r�T�?:�;���A��#�P:\����u)�QX^�2���@i"M6f��������5��	"	���?��o��N�1�a�g��ۓyP������1��
O?�p٫j��"�yL�x���Ys�}�q��?Xٵ��5�,����F]�J�������	UQQ*rb�5��6��uF�p�	_�P塙@:/!M_[V�I'�
n� 70^�d�e»�-0^��,�:�	S�uP�M�zK!�g٪�'�)��F�p�	_ى�#�9�$�oWU� ����L�m�C��#��;����B�	?�gwC�N�O�lK���K)��F��P������_#Ǚ��R�����'c.�	?0-� ����Jv���,����@p~�@oH��{T��qɮ����D���,%GJ�=�rW�K�v��|�5������zWG����ʙD�0@]�����>'�6�*�q�t������ϩU�R�4�t������:Wp<!���I��d�>�r=D�9�)�Ί#|�Ӏm��!Q	s>R=��@�wG�ɽ�&���[�O�VG/"���@V��"W���à\j����f���ԝh<K��}|�?�M��\%i�������E�!��o�8���RX<���O��"P)�6�m�`�� P����Y6Z����*y����,��/�&�5K}�*���ՙ��e'�������s�SŠ��z��Qd_No���?�%6=�wۛփ��A���ƍ�sv�{d�� h�����\4�뤯r�J?Ȑ�����Bbp^�ߣ�y+dꜱ+�	Q>���ě�T�t�g��W먎�E؝,}����bq f�&�������1���?�~ .��ԟ����A(B�������%�R#l���[�R��0)I�P�z\er�G������t=X��Q�k��/�m�K�֩XQ0)I�P�z\er�G������t=X��Q�k��/�aa?\��E�h�,�B�Q�#K
�SI0��<҂�H��T}t%:3VU=f�:>5��Oh`B�VT�́B��h�G#o��c��Q�w�)3��Z�����ū=ċ)$����W<:K��{v����<�OF�P�]�Ҽ�w	�I�D�J�Vc���d��x�OB$��~��WRKD�vQF'�BI��^{g����M�b�K1�>�yl2����ar��Z�.��n���=�W�^a��	Wb�tm�5��Oh`B�VT�́b!���J�TҘ��S��!�`ڹ�m��!���~��WRKD�vQF7��� h)��Rd�'�U���'����\�<�f���t��F z_.?�P��Y��G�y	J�X쟋�yN�F�8I���W<:KRKD�vQF'���_<+��c��k�:���"���0�g�Qt���~��WϘ���F,%a�(#'�4H�KV��iI�yl2����ar��Z�.f3���W��J�9��E�M��1����{T�_0��ݤp\�Ì��I>/�4	���] ��2��wt�,g� g�Qt���~��WRKD�vQF���<����(�4#ᓠh�A�f���� ��#*����Z`ύ���#���WdꨞR�"�/y������9:F(H��u�6�S��}DFB�5��M���>���6����_��l�ֹ�TC�r4��%z�r�sb���t�V/����!D.-#�L��"=I��`�^/������N�������ZMӼR��F}��d��3ic��ݤ�����a3m �)\IEs�1��)Z؋$��,!����9���7,���)D����U����H�;��A�YyB=�u�@3C�����շ���=�Z��K�`؋$��,!����9��ɽ�*<e�˵�L�2i5b]���j��x�3KuJ:p@مI���?�G�Y?�FA6����L��Թ��<G���"��+�~��ԧ$���i�'�2�5��Oh`������<嶡+U�n)�&�|�D����L!T�~7 ��!Jx���]L�E�����I��嶡+U�n)ɽ�*<e��s2�E;N�lU�+�+�1��@f�����p��}�tؤ�l�k���,(n0�Q{�5���3��z5�g>X���rt?g=T�`N=L��,aM��5��<ɽ�*<e�];�ٻ!Ŷ�,�k[�u:׈S�y|��5�L/%�QH�#D=[�����J���C>��M �V��{u�8I�f]U�S�#��˥ҳv��!/�n�]��CH�v��
�YX�#�y���dk>��E�qi/.�ͼ��ow��"KB/�Z�0P�+
$Q9sNy��n����e��{�KG��u�`r�_Y�o婛�F��K�G:�]v�`��Zݪ+il�.SM	B"�3��[$���J�m�p�id��H p~�vo	u6��������~Mv��*��W�+�g���Qt�%��٩���W&���}��]]W�k69O��=��7���l陯�'¢c*���lnr�����5��?��Ͽ��~^-C;xc&z�j��S�#��GEW6�7@-o��:Q=c@�LT!���O�0��͍��aK��N�ow����u���5	v�aH���&q���g�i�r�rz��F��$>@77�D^�]x\��斳9��u�h��
[JJ����W<���Na��<��g��k����k"�Y���ߢ?a�\OW���<x
����s���é;�Z������Q޶gqw]V�ȣU��;:�=�EBi�G�"�e���#�S0�zdr��#��m(�D�t26�U�ئ7�����;���/Ty����jc'��/(JO��K�^�4�d��=OĪ7I�\�v��⢻��d~�}sC�q�=�TG�����Y[v�_�8���1��$��u��}y����B�]3�#ս��F-��m��@�-��/�e��L�gB ��2A�v)̻y\��TUɇ�6������)�wi�n �w�ny�2�d �|w�Q΀�zSD�X�a��њ�0h�����G#\�0�����Ӆ��%���8���t���+�W�D�j��P�FK�M�z���}�C������b���K�e�1���|"ÝWj:�,��Y[v�_�BD��Kũ�V=z�iwHm�H��7(+�˹��Q��B��]��_�L�fp���(�HS|��(߀Ď�\b���Ori ,�顫v��,5/���J� @A�˘+�)������^�]�X���:Ҽ.�:7�!�P1s$�8�W��x\��斳.a�%8A�V$�__�;�gV=���,3��n����˲|���V�X�z���sO+��RYc�=$�[��x9�G�S�#��x~���`�7��{%Ĭ��'l�X�.x\��斳���J��^o��fy�]ÌJ��,�J;xc&z�j��S�#��F~Z'�Z������H�ayL\�3刅x\��斳���J��^o�������D����២x �t�6\�3!PƲ��uMG�
H ��E,��RK�"�-��H p~�vo	u6���^��:�|\���}��F-u9{0��%�Zݪ+i_�)�zy�Bwfax��M�2������]x\��斳���J��^o����Nހ�kx�<.h��@*��wl6-��Lv�fJz�"4g~K8�9`oM�r³t����2I�յ*s*���  Ƚ4n��G��2�dH,��\����2I���-��&��?�/�oCG��=%K�eIi%$����J�P�u�{	}�g�:~�N.t���y�P��{v���ɉ6$�獎\�v�����Z�k�5�*N�s���E9�)�V'�s�1FT^�L�����2I��v��x9�Bs�]��b��_��i%$�����֍5\�+�Ayɲv$Y�vN�rt���y�PU���ئK�}r!b&X͸8yw�T��Fz: ����^-��8"���)��DP.�'�@k�{��������L�8jɽ�*<eb��_��i%$����J�P�u���9-�m�\�-�k�<��Š����ɽ�*<eM)���Mz��]'E���id��H���Hi޲39���H9R0|c���=r���4GHt���y�P���qE���	+���e��Wx�����G��iP��[P���<Q,�X�Mة�ՙ{�4}���Zf�O7H����HO�F]�{�ɽ�*<e���Z�k�5�*N�s[�%��+�"�ٓ��	G�-�k�<��Š�������g)Y+�_xZ��C���~�	N�.X'.86|B&	���o���͖����E�T^�L�����2I��9��w��1�*ݚs���E��ɲ&st���nđʘ�F�,O��gߋ��-��8"��-d�4)���ɲ&s����P����<Q,�X�Mة3�9�D�Zoa-�[Ƭ�WB�W�����|��$���]�L#-Դ���V�>H��yz�3?��V� R�T��k�X�~{+�	���v�dq�LU�W�X�Mة�W���ZB�:��n{%�UdmB7 ���Zm�k.\�&eu����>d$q��s�C#e�u���g_���P�`��՗Έ4LkFl�Ym��#z�L�D,)�U���~��.mz���D*˵q%��A)�^U��[�f���y���b�g�}����u:?̘�3#;j��=�`��Έ4LkF�=�r|�Hi޲39���H9ӁbF�i� ]�ʺ����Q�X�zι�@�[�M.�r�Ϫ9��P�	 L���`�1�:Nw��Ҩ5$�)iA6���^/a�1: �18e���zG>d$q�	�덮�pO�U���~��:Nw��Ҩ��>���*%��8Y]���(�[�v��,�b�FhwI7Is[���ɽ�*<e�LG��3�\0��;�O��ӁbF�r����i�'�]'E���i���j����t�(v��T^�L�����2I��Iu������O����`�v�P�5� R�T��'8L��t�q\'��=\�
?��"���<Q,�X�Mة��_QSżtX�zι�@�)K��g��T^�L�����2I����zbZ�9Hi޲39�)K��g��M)���Mz�E��7ۅ��ycxB}��ɫM�����2����5c	�s~;fTE��7ۅ��&ꬶ�R�M�����2����5c	� b��N�
�I���Z������6��5�hJB�G#y��I>/�4	8'�"7��lT�:��	����1C��uԅsE%��D�&��ö�#5��{v����<�ܥ� �R�ߴt�D{�h��@�ɵ��g���>���|��[����;t�����	�~��Sx�,y��ש�zk��b��M&���Z�k�N�ʆQ'�H�e�9V�$�S�g�-���3���T..+`��M)���Mz��?�Vl��n�b>L�M��pRV���ޡI���W�Y��xlYE��7ۅ��&ꬶ�R����4���j1;�J�Mc(J ���"��m�
9Gi
��Cj�%�u�){Kt.�댴]�S�g�-�I�2��eo��H�>��.��^/a�<!!�DIB���a��{e�cŬ�W��w�g�˴�m�3'k:�<�WV
v������Q��z�`u�t�W�/����K��'K�{�a�.��U&ځ"�*	�}����u|����x.�R�ߴt�D{��ש�zk:��|��;�Y��##����?5�J����<�`��g�ḋ3���Tf�2N�2��}!�Lڜ��[��L�)�>��X�g�U���9�iP��[PT^�L�����2I��3̧牊I�eC�O�|ˎ�D�cyHt���y�P17J m-Q�~�LZ�BJ�bZJ{�[��(`�*���r�i1��1�C�j ߥ}t�6�&���pO���~"������]��f�1��e��M,����6�w��dg;�f�Y��^/a�Hn����y�֠���ɐ6]��>�����E��7ۅ����zKa�PI�$NZnx�5�{}����]C	à�{v����Y5V���@<�$���ɲ&s����P� �E��7ۅ����zKa�PI�$NZnx
9�������I{'��+�_	��������FL��.����J�^����'�����2��z'��x}���{H�3���.e���D�f`KK�Î��w_F2]�J8���@�q��F2]�J8��X�����cF2]�J8�F2]�J8�	xG}�a:����"'2�I� ��K��w'ä
_[FBQ#�dtt�q��Q���p49�1��g����b���rM�׻�m�Î��w_F2]�J8���@�q��F2]�J8��X�����cF2]�J8�F2]�J8�	xG}�a:����"'#d���^d��w������M�D8U"�����aZ7P��/���	MU%^"-� M�׻�m����M�ؾᯰ����G�J��D��:������Oz>+u�N*�麁�9�#/M�=C�\:����"'#d���^��7�ٚ*���M`�'��거���aZ7P�k_fè�s���K��uM�׻�m����MG��{$�'����G�J��UJ��ٖ�����Ozɽ�*<e��{��M�=C�\:����"'<����u��}/��<��P���M�?Q���aZ7P���G���Jδ_��uT�M�׻�m�Î��w_F2]�J8���@�q��F2]�J8��X�����cF2]�J8�F2]�J8�8DR*�h�эYR�w1�$�q�H� �!�bON)�5eĊۏ!����\[/��_�].?� <�����\��4\�g~18�3�^�2hZj����-{����>�ko�U�����q�!��	m���3� �`Y,�R�׉��A��Q����_��Tݥ/��jma�WY�g�L������o��Ϟ�	���Q���n�Ѱ�*}��Pj�$NZnx
9�������I{'��+�{�R�I#-Դ�� �`Y,��S��A�8V�al�[]$5��hޅ����/H#-Դ������_*�YZ͆ˎ�V���5v3UF2]�J8�tQٍ��^F2]�J8�tQٍ��^F2]�J8�F2]�J8�F2]�J8�wԧ� �n:m5�1g$���Q����HER�M���X֖����)P@�zz4���_I�ab���b���r�"� �
��Y{��6X���l��D��	���e���^E��s��/��7rٺ'њ���I{'��+��n�<�ӂ�ѱ~C�F2]�J8�ƿ�bqF2]�J8�ƿ�bqF2]�J8�F2]�J8�F2]�J8��Se�����+/r���/�ᢤ�ɽ�*<eۻ���T�'ɽ�*<eu���(+䩾��k����~�.>��M�=C�\:����"'#d���^4`!������ۉ�J���ɽ�*<e���M���Y��z��/dx���������ϖ���8��C��4�L]�����$����uc;���7�ٚ*	?Kʩ�䉒CD��< ��+��z!�JE���D���*���ɽ�*<e���5��8P?Ω�����DhY��F�쐠�g��	_��k,�>7Y�����5�T��I/YZ͆ˎ�u���(+�v���N�Ax������|	r�x����/�ᢤ��t�q.U���}^�ć�M�׻�m����Mv&�v������G�J�F.���щ���G�J#d���^� �c]�4�����L�L�"� �
�[��y��3`� bL�d�������Oz/�v��ER������Oz�C��4�L}�"�:H�{Sڥ�W,��������*��?d�3���X&*�Q� ���K�����N�s��Mi�R�ɽ�*<eFZ���m�ɽ�*<e�P8񒽮�ǅJ�nF2]�J8�F2]�J8�V���5v3UF2]�J8�V���5v3UF2]�J8�F2]�J8�8DR*�h���A)�^U���H��8ܟ��Dz��JN*�R���D�m `���*`(�l�pۨm�4j�N�
�I����c#��~�����Wdꨞ�E��Ee�l��h�*���Z��������v�j��tc�XF�?��.���l��o+m�غP��`�a�5,�-8�Y�&�9\�&��X��f�֗۬���-�.�t���%D�M�V��Ŀ�>J�g__�4D^��_��b��Z�p�+�n�/�G��Q�֡�$���cW΀��˺�1��?k��$����cW�Q��z/M����v�j��tq���g�� ��Ԫ�N��+�� �z*B���C;}�J���WW�iw3A�ώ1�Đ���A�8.h�,1z|��@|=W�������~Mv��*��;���s&��%���PlS�����*��Z²ǎ�U�#�.����p��y�MWO���5���@Ԁ�r_�g-���gLٗ>�^�p���[#�����-��6����eC�O�|ˎ���V�uCM^��D�}K-��6����eC�O�|ˎ;}�J���WW�iw3A�ώ1�Đ���A�8.h�,1z|��@|=W�������~Mv��*��;����n������PlS����`���$���
?�	���3�T�JS=�ҋ\�d��	_�������p����;?Q3�0��J����p����&Z��&�K�z#.��(�;�")8�^,3��0ddRy��5��t�I:���Wdꨞ�E��Ee�l�kI��ϕU9���
0U2ZF���f^��_��`�ր������bo8�Y�`Dn�2j���N�o�VF�NŐ!}�&���pO���~"�Dr9V�Lʇ��t�isCܛJf,�1��d�ߪ�q�7�eC�O�|ˎ���V�uCMU��`���5����X�*�^e����1AiD���cW�rr��!U��NV�q�.��Ԫ�N��+�� �z�*�^e�+#�r�5h�kI��ϕ���d��X�;��μ��M��)�Q�o3�� ~�������DLc�w����'.�v�a9��	���Ǖ[���I�%�c������Q�M��䕗��v�j��tc�XF�?�7�gv;&��`V�f�Bɽ�*<e���+��ͮ�F�ģ�M�3pI^C�����p���q�И�mJ��E|�m;ɽ�*<e���<���*B���C�H
E#LPA�Y��g����,�4�
�9����j`▘9�U�����@�P�=�����P�OP<^�e}Mmnk���,(n���<����(�4#ᓠ���H8��s�[r�/���P�OP<���A�]�AX슚Φ_o��u�삙��q�E�Sga�������<�<�XS�<)�	H�e�9V�$�S�g�-���3���T�X"��|���@z�J����@��K��'K��HL#-ׅ,�g'P��S���=,���V��9�p�پ� �+���Xw�gR��{�g��(e��>���LC0%�Y[v�_��~��^��R��\�P�6�J�KD�/���z��ɽ�*<eu.(�B�3d��pl�R/A�}QW�Զ݈�}A�����n��rɽ�*<eV���5v3U��@�q��F2]�J8�M�F܅ڀF2]�J8�tQٍ��^��@�q��F2]�J8�Ƣ�����x�\�u/!����֌�����ku`}�� �@Rf�=�Rt�-z��rٺ'њ��I�����*D�d�ka|w�kK��%�w�8Y[v�_�����@JF2]�J8��#�:�>ƿ�bqF2]�J8�F2]�J8�%w�
�H=�#�:�>F2]�J8���o�s��NM{9q��F�L$������3FcgGqT�&g�b�Z���wk�{�|o`����mX�n\L�l߲!w����@��ǂ�VJUT���)!)gP\�L���D�)��R�S����
�L����j�pSQɽ�*<e=@�����W�^a��9DcI���JПE�[5ɽ�*<e��
����)�''�!h�X�>�z��`V�f�Bɽ�*<eɽ�*<eJ/x��8�4.Ee�T�����^�^Wދb	tɽ�*<e'$��R��eL�"۠��JПE�[5ɽ�*<eɽ�*<e��`V�;�.
����d�x~���`�7��|�Q�ɽ�*<eP�7ٝGy�ɽ�*<eɽ�*<e��Q��mD�m��nN��o"/d�m��k �u+�%0ɽ�*<e�´Z�zY+{�G%��NIL��|6kcb7A�Y��gɽ�*<e��JU׶�7��y��� TO���A�:Nw��Ҩ����p��ɽ�*<e���Zf�O7H����H�NIL�h�Ǳ��mɽ�*<e,4���?w�0���=�Hi޲39���H9�^.|�M7ɽ�*<e�����>��ɲ&s�-�k�<�GaX-!���NSad��ɽ�*<eF#���	��ǵ��������r� ����[Y�ɽ�*<e?tB��XT�S����Q�^>v��(y����]�������� ���B;ɽ�*<e�J�!/�:��n{%!�׃>8��NSad��ɽ�*<e����Yڤ	���v�d��
�0�_xZ��C�ɽ�*<e��ky�-��|��������i<�R{E�6��h#A�Y��gɽ�*<e:`��r�rٺ'њ���I{'��+��CqwɂjO�F]�{��E��-ɽ�*<e�
�9����ɽ�*<e��P^}Q���S#��\[-�H���Gޛfe�^C�ɽ�*<eɽ�*<e�Q��
ձXt�G�
co�]+nO�BT�\�V��Ԧ���=��a�h��~z�j�=��=ɽ�*<e,4���?wɽ�*<e����Ʀ�ɽ�*<e�oc;�Eǎɽ�*<e�)��8y�����p��ɽ�*<e�ǅJ�nF2]�J8�F2]�J8�V���5v3UF2]�J8��#�:�>F2]�J8�c'
fg��rɽ�*<e����8�rٺ'њ���I{'��+�ȵ�m��O&V�Zɢ6�%3�VA^����'�r�#��"�ɽ�*<e����n��rV���5v3UF2]�J8�tQٍ��^F2]�J8�ƿ�bqF2]�J8�&MQg��/Qɽ�*<e�VJUT���?�(<��ɽ�*<eS���u:i�i�r��qi��ߔG�=��ɽ�*<e@�^�~=fJz�"4g~֖�9���Iɽ�*<eɽ�*<ex~���`�7-�a�(%-U������ɽ�*<eɽ�*<e�o|6���I*<�����Y���锸��j Gɽ�*<eɽ�*<e�´Z�zY+{�G%��NIL���a��C&�-�k�<�Fb�9J��90H��r�dZɽ�*<eɽ�*<eO�
�����=��"V�wo"/d�m���O05�j��ޛfe�^C�ɽ�*<eɽ�*<eɽ�*<e0����� ۄ�v����esȜX5	�l�khy�ɽ�*<eɽ�*<eɽ�*<e1��0ɽ�*<eɽ�*<e1��0ɽ�*<eɽ�*<e� �O_¼��"�	� �3�\0�k��6uQ��xLj���S1��L�ɽ�*<eɽ�*<ey�?Y:�B!�]�Z'�x���]L�Eɽ�*<eɽ�*<e����n��r"*c4Q��e �Sծ�=�B���.���X�ɽ�*<eɽ�*<e�VJUT�����B��I!U	��+*���{�ɽ�*<eɽ�*<e�'1�*��P�K��_�t��>^��%$��x��%>��^���	�ɽ�*<eɽ�*<e���R�n�eN�:�$,=���G���y�w�c̗��Q~�Z:�^��.�Ȉ	XC
�V[�ɽ�*<eɽ�*<en�{��G�P�K�Ҁ-�k�<� �y1�P���B���������p��ɽ�*<eɽ�*<e.\��O۳�xLj��bWk؏э0+l�.��O����`3�s��Y�yO$�,�ceɽ�*<eɽ�*<e�p\�Ì�^����'V��Pf���$�>�P��v�.?�}$/Xp��ɽ�*<eɽ�*<eɽ�*<e�`�����z�'�|\�/J
��r�L	�n_ɽ�*<eɽ�*<eɽ�*<eʛ*~�9N*@o�JY�H
E#LPA�Y��gɽ�*<eɽ�*<e����,�4ɽ�*<eɽ�*<e����,�4ɽ�*<eɽ�*<eh�p]h	���su,Z2�Hi޲39�)K��g������p��ɽ�*<eB1U���vܪ0�:pHkn�f��H�ɽ�*<eɽ�*<eɽ�*<e� �O_¼���f"k�<D>������ɽ�*<eɽ�*<eɽ�*<e�O����`����+L�
��-R�DŞ(4������JrAɽ�*<eɽ�*<e��Lm�$�o̗��Q~�Z:�^��<�b�A���H�w`l�o"/d�m��.��l �rɳ'ԙɽ�*<eɽ�*<e�پ� �+��7�]O�#-Դ����c:�_���*"�̩(2N�uV�:�ɽ�*<eɽ�*<e����@��
�늎��	���v�dj�?m��������ɽ�*<eɽ�*<ex�m���`�υI��psZ�跐UW��@z�Jɽ�*<eɽ�*<eɽ�*<eN5G �):B)�[f3��`��e�d9Y@��ɽ�*<eɽ�*<eɽ�*<e���M��#-Դ�� �`Y,��z���}�ޛfe�^C�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eX�zι�@�}�V1����P�,&f0H��r�dZɽ�*<eɽ�*<eɽ�*<e�+�r��y�ɽ�*<eɽ�*<eɽ�*<e�h4�+�t�q\'�������C�oCƞ�Xܳ��_�2�ɽ�*<eɽ�*<efD@t�u��䍀�<��Cqwɂj�NILș���!BM�c|���	9�U[j�xOɽ�*<eɽ�*<e'$��R��e�����kV�ɽ�*<eɽ�*<en�{��G�P�K�Ҁ-�k�<� �y1�P��1l�XiI�����p��ɽ�*<eɽ�*<e��݇%����3��H�I��0+l�.��O����`3�s��Y�yO$�,�ceɽ�*<eɽ�*<e"7�!ne*5�L�x;��@�֢ޮ�H,�a��(-y~�I}� ɽ�*<eɽ�*<eɽ�*<eʛ*~�9
���"��H
E#LPA�Y��gɽ�*<eɽ�*<e����,�4ɽ�*<eɽ�*<e����,�4ɽ�*<eɽ�*<eh�p]h	�E���l�sfHT�N�g�o���S��hɽ�*<eɽ�*<e�`{�H7��ӯ�oM�k��3'������p��ɽ�*<eɽ�*<etʐ�&'���Gq��s]�j��rM�#������ɽ�*<eɽ�*<eΡ���8�u�$�k ����ԥ�X�U2�f$�xKɽ�*<eɽ�*<eɽ�*<eM�L�uP�@����?��Q����2l=�ɽ�*<eɽ�*<e��}Gδ�-��x�f�Up��	f��"�`V�f�Bɽ�*<eɽ�*<eɽ�*<e����Yڤ	���v�d��
�0�_xZ��C�ɽ�*<eɽ�*<eɽ�*<e�[U��n)*ݚs���E��ɲ&st���nđʘ�F�,OkVib�(�`ɽ�*<eɽ�*<eɽ�*<e0��l��hHi޲39�)K��g��ھi��͗
ɽ�*<eɽ�*<eɽ�*<e;O���Tu�� ���I~W���
���aˉ�rR���	?�Z���L�8j�dY)���E���I稚Sv�K{|T	���-�8wɽ�*<eɽ�*<eɽ�*<e�����K�B)P�B�*ݚs���E��ɲ&st���nđʘ�F�,OGaX-!��t���y�Pɽ�*<eɽ�*<eɽ�*<eAjC����?At�#�<��a��X���l'�{�z���ƾ��e湘��� � @<�$���ɲ&s����P� �����p��ɽ�*<eɽ�*<e��8t��6nh�
nɽ�*<eɽ�*<e��8t������p��ɽ�*<eɽ�*<e�ɜO �H70tW%m����L�8j�Or6u�m�e��Wx�����G���d��+RA�Y��gɽ�*<eɽ�*<e��`V�;�.L�&�$��:$�m״HT�N�g����3�86|B&	���o����f"z�7�~���#hɽ�*<eɽ�*<e���(���"�&��&P�	G�5�3i0�,|gW���0}B�ɽ�*<eɽ�*<eɽ�*<e����X-�9;j��=�`��Έ4LkFRu�d�lHi޲39���/�F�`V�f�Bɽ�*<eɽ�*<eɽ�*<e<vy%�p0p~W���
���aˉ�rR���	?�Z���L�8j�j�J��~W���
���aˉ�rR���	?�Z���L�8jGY��J�hɽ�*<eɽ�*<eɽ�*<e�<�ܥ� ����,מ
��	�y{I�7�P�,&f0H��r�dZɽ�*<eɽ�*<eɽ�*<e�э�&���;���8���^p�!PU���[��ӳr���?��t׉s7�yO$�,�ceɽ�*<eɽ�*<ef�{��t�ɽ�*<eɽ�*<ef�{��t�ɽ�*<e'$��R��e��Ω-b�ɽ�*<e�v��,��ɽ�*<e9�ݞR��=����n��r�\�Zai�����wD�N�jێ�ߔG�=��NM{9q���z���^Bɽ�*<ea�_��)5��㬟S/��V!��:^��J"�VJUT���;E� �21F2]�J8�tQٍ��^F2]�J8�V���5v3U��@�q���CMNY�ɽ�*<e��Ӿ�����D��b�~�	8�[��+�r_�j�T�U�/L�י(KC�Ɛ��$7۹Xmɽ�*<eӂ�ѱ~C�F2]�J8���@�q��F2]�J8�M�F܅ڀ�X�����cƿ�bq����p�����/�rQv�ϗ�1<�k�:HW�?��s�G�
��2Q�W�l��R�ӫ�
���"K��b.����p�����HG��}Gδ�-��(ʂ���<��"֧XS�<)�	ɽ�*<e��9V�N��TҘ��SJBD��m�`.苢��w�ɽ�*<eɽ�*<e����!~p�֢ޮ�Hy����~����p��ɽ�*<eU��a�>��J��Y����.����l���G�J¾al�%g��4PH�Y2�hv����D���dQ�h�͝ɽ�*<e,4���?w��cϖ��L8��\Ŭ��G����_�2�ɽ�*<e�{o����T"#��rxB 5�yc������ɽ�*<eS�/Y:n|��U���~��:Nw��Ҩ���H�h��Sz�̞��ƒ1*8"Z�d0H��r�dZɽ�*<eɽ�*<e������ko"/d�m��{-�[�WUIG=M�؞A�Y��gɽ�*<er�֏��9��W8 �+N�����p��ɽ�*<es�5�|Y��{��������L�8jySۨ�P��n���@��yO$�,�ceɽ�*<ef�{��t�ɽ�*<e�VJUT���51=�(��A��-�N�e~�5���qd�ơ�ɽ�*<e�'1�*�|�JnQo1l��`ؠ���x5������8�!�|ɽ�*<e#�^�����	��ovP�`����Z:�^��[��M3)�$ɽ�*<eۓ]d������`�1�:Nw��Ҩ�E��o��ɽ�*<e�VJUT���h����Ny-���qoYy�֠�㙳���,�+�duX�O-��_�2�ɽ�*<eΡ���8{��<訄��j��p_E�)\�?�.+:*CgI�W�#$ɽ�*<e�i{ޝ��i#-Դ���X"��|��R¡�ɽ�*<e���Ɔ��"ɽ�*<e��9V�N��TҘ��S\��b&gLB�`V�f�Bɽ�*<e�VJUT���?�(<��ɽ�*<e��d6����ɽ�*<eɽ�*<e]~�����ɽ�*<eɽ�*<eӂ�ѱ~C�F2]�J8�F2]�J8�F2]�J8�ƿ�bqF2]�J8�F2]�J8���o�s��ɽ�*<e:����"'ɽ�*<e7��� h̚Ff�(#�ɽ�*<eU��O�ay�֠��}i�?ܻ!ɽ�*<e?/8V7�&�F2]�J8�F2]�J8�F2]�J8�F2]�J8��#�:�>F2]�J8�	xG}�aɽ�*<e,4���?wɽ�*<eɽ�*<eRr�t5��JmP��8��IM=Cfɽ�*<e��ʧ �e�>*�����ySۨ�P���&-�����ӊ$]���JrAɽ�*<e7�ϙ��&'<|f�z+�SWĞ�ɽ�*<eɽ�*<eaL`<��x�{��Y/���z'��x}��u�^�d�X�zι�@�)K��g������p��ɽ�*<eB1U���v���`=��JПE�[5ɽ�*<eɽ�*<e��F�#���ٓ��	G�-�k�<�GaX-!����-�N�e~�5���&�K>Z����-�8wɽ�*<eɽ�*<e�VJUT����C��4h��:M�&�m�Z�YK_��L���J�ƃ��r`�>MFD']4`G:G{�"Y�TndX!(P�|na��+����p��ɽ�*<eɽ�*<eB��iA����E����o"/d�m��N�z�eo>tޛfe�^C�ɽ�*<eɽ�*<eɽ�*<e��}Gδ�-��K\��)�Z:�^��f��*%�)c�`V�f�Bɽ�*<eɽ�*<eɽ�*<e����@��K��'K��HL#-ׅ,�g'P��S�,���~N�'ʆ�%jȆ�)���A�Y��gɽ�*<eɽ�*<eu:׈S�y|��5�L/%ɽ�*<eɽ�*<e����,�4ɽ�*<eɽ�*<e��
���Դ��M8�M$TrU:Nw��Ҩ�s)|����x���]L�Eɽ�*<eɽ�*<eɽ�*<e�cG�^k�{��������L�8j7�j�!�k���,(nɽ�*<eɽ�*<eɽ�*<e��ky�-��4.Ee�T��T�y%f�v�� ?ɽ�*<eɽ�*<eɽ�*<eɽ�*<eX�zι�@����7ě��w`&�j��:��P�?#����������z86|B&	���o����N阈7�>	D�k�<�a��xLj�������w/rA�Y��gɽ�*<eɽ�*<eɽ�*<eΡ���8{��<�Tϱ'���W��<iVF4RZ�utk7��K��'K��HL#-ׅ,E�����2=�4d3A�Y��gɽ�*<eɽ�*<eu:׈S�y��L��Ԝ�x���]L�Eɽ�*<eɽ�*<eɽ�*<e.\��O����+kȵ�LE����O���E�ɽ�*<eɽ�*<eɽ�*<eS�/Y:n|��U���~��:Nw��ҨƮ���0�v����T��&�K>Z����-�8wɽ�*<eɽ�*<eɽ�*<e����@��K��'K��HL#-ׅ,�g'P��S���=,����NSad��ɽ�*<eɽ�*<eɽ�*<ef&L6��ĩ%�<(���Q�����p��ɽ�*<eɽ�*<e��8t������p��ɽ�*<eɽ�*<e�+�r��y�ɽ�*<eɽ�*<e�+�r��y�ɽ�*<eɽ�*<e�����E�J���O������ɽ�*<eɽ�*<e�'98t�'�-�k�<�GaX-!����K\��)�Z:�^��.�Ȉ	XC
�V[�ɽ�*<eɽ�*<e#���-@f8��\Ÿ��M2x)M��ks��JПE�[5ɽ�*<eɽ�*<eɽ�*<e�!B��'�Z۰�E>wGg	 �'��"���3�-�&ea�k �u+�%0ɽ�*<eɽ�*<eɽ�*<e?�/�oCG�V��\��?�6pΑĘ�ɽ�*<eɽ�*<eu:׈S�y|��5�L/%ɽ�*<eɽ�*<e�ٍ�t��OiҢ@���U*��	e �J���v7�7ͮ�WчP��kt#��=7���6�{�XcN��o��Uj�D�;����p��ɽ�*<eɽ�*<e�cG�^k�{��������L�8j�oM���4k���,(nɽ�*<eɽ�*<eɽ�*<e�M��������6Ɯ�N.8��l��:4�GN#-Դ���V�>H��y��`�7.\�ɽ�*<eɽ�*<ef�{��t�ɽ�*<eɽ�*<e����@�������=�zt(xw�mӁbF��f����ܮ���ۉ+?�_1���e7z�]�rY��c��H��U���~��:Nw��Ҩj.��~�U���~��.mz���0��ɽ�*<eɽ�*<eɽ�*<eۓ]d����
����d���'#�H_hʖ_�*(�ɽ�*<eɽ�*<eɽ�*<eۓ]d����L�&�$a�\�Y#-Դ���V�>H��y�¼�B����䍀�<��Cqwɂjp��\�;$K�/��7X�zι�@�)K��g�۫[jj�ɽ�*<eɽ�*<eɽ�*<eӳr���?�t�V�,�X�zι�@�}�V1���&����sj��.��cۘî���^ţ�U����S�+hO����p��ɽ�*<eɽ�*<e�+�r��y�ɽ�*<eɽ�*<e�+�r��y�ɽ�*<eɽ�*<e��'#�H_h��wt;*!x���]L�Eɽ�*<eɽ�*<e.\��O�P�`����Z:�^��\>-��#-Դ��o"/d�m��.��l �rɳ'ԙɽ�*<eɽ�*<e/�e�=~���PB��+6L�j$7�-�%E�}��kx�\B�\1{�E�@E��V�Z&eu����>d$q��6���ɽ�*<eɽ�*<e3ƹq�nNs�ab���-�k�<� �y1�P��Hi�Yex�����p��ɽ�*<eɽ�*<e����n��r�#N�K�$,����^���+�a��{�)(�X����*M�ʐ��&ѩ�&�Ii���m�'�EA��[/�����x�ETOf�25����p��ɽ�*<eɽ�*<e����n��r�hn�@�L3�|C�@D�K��'K��ǉ��������� ����t@BA �粭�@7ָi�Z$ݜ?�9��7oa-�[Ƭ�
��,�fM�ɽ�*<eɽ�*<e����@��K��'K��HL#-ׅ,�g'P��S'D�v���.gW:?�g,�&U���Ϣ�5�RM��R��k9��:;��2��:7ɽ�*<eɽ�*<eu:׈S�y|��5�L/%ɽ�*<eɽ�*<e���M��#-Դ��Xi�q����_�A�����k���,(nɽ�*<eɽ�*<eɽ�*<e�� Z o��޿�ة�V.gW:?�g,XFC�6��Nqb;e�Y;t�q\'�������C�oCƞ�Xܳ��_�2�ɽ�*<eɽ�*<e��
���k�}�1�ع_��`�����j;�����p��ɽ�*<eɽ�*<eɽ�*<et�q\'�������C�oCƞ�Xܳ3�>�Z�=5�3�\0��;�O���yy�=����
:��{gɽ�*<eɽ�*<eɽ�*<e����,�4ɽ�*<eɽ�*<eɽ�*<eZ��#1�oa-�[Ƭ�ƥ,`��u�'ʆ�%jȆ�)���r0+�3���3�\0��;�O��h����=1z4���_I�ab����o~S~�[��A�ɽ�*<eɽ�*<eɽ�*<e�[U��n)Ꞿ�?�tS�8���j�)���F��> N
��ز��'^0dSQ�L>��ƙ)(�X���n�x!��4�k���G�����ɽ�*<eɽ�*<eɽ�*<eӳr���?�t�V�,�(�k�>��D�ծe�o�U5Hv���"���m�j��.��cۘî���^ţ�U����S�+hO����p��ɽ�*<eɽ�*<e�+�r��y�ɽ�*<eɽ�*<e�+�r��y�ɽ�*<e��8t��^�$`#^gɽ�*<e�
�9����'$��R��e�_o��u��p4�8��m?�\�v����(��H�O�
����Y�x=�U�#5����F���c�H������ �
����ܤM�Yr2�(���<i��=����/�žCɽ�*<eZ��z}L�|Ǌ6��[����m���s���9�� �+�`�Pɽ�*<e�+�r��y�ɽ�*<e=@�����W�^a��P�쑱�JПE�[5ɽ�*<e,4���?wT�=P�������o�*͗�O���ɽ�*<eZ��z}L�|Ǌ6��[���.����;�ɽ�*<ef�{��t�'$��R��e�_o��u���پ� �+�S�&,dNgƧ)����L���D�)��R�S�����I�%m}5Ek���,(nɽ�*<e�~l��.C{g����M3i�!��[�x���]L�Eɽ�*<ec�t��]�,�U�n��K�c��q$�(�hY��aȩO.�����P�OP<���A�]��[�T���e�4Z�[��lc��hp�{b!ɽ�*<ef�{��t�ɽ�*<e��P^}Q���S#��\[-�H���Gޛfe�^C�ɽ�*<eɽ�*<e� �O_¼
^��qυ�A)U>6�a?ɽ�*<e�c�!7�Ch��iv�������b����Ȼ:Y>�9�JY���$��w�?�PÂ��(�ɽ�*<ef�{��t�ɽ�*<e��P^}Q���S#��\�VV�*H�ޛfe�^C�ɽ�*<eɽ�*<e��H��8܎�$���������N�t���y�Pɽ�*<e�q�И�mJ��E|�m;ɽ�*<eɽ�*<e��H��8܎�$���������N�0H��r�dZɽ�*<e�+�r��y���8t���ߔG�=��{��/>�d��i�M�.����@����+�(G_�x���ޛfe�^C�ɽ�*<e��}Gδ�-n;��w ����7U��p������p��ɽ�*<e,붏�#�|촣�yOK8�j�=��"�NR�j?ز�<}��V����F8��1g�t��ڭ�b�o/�n�]��F;�d(���_%lɽ�*<e����,�4ɽ�*<e��9V�N��TҘ��S\��b&gLB�`V�f�Bɽ�*<e�VJUT�����B���LI�${�ɽ�*<eɽ�*<e�Bs�]��ySۨ�P��E����'{���of ���Zn���cь�+�`�i�]Kɽ�*<e1��0P�7ٝGy�����p����;g`��I6P�V�����p��E)z\ː�ԝ���a�pp9��jx���]L�Eɽ�*<e=@�����W�^a��9DcI���JПE�[5ɽ�*<e���a_��{X�aҥ��!��Y�N:��6C�p����P�ɽ�*<e����,�4ɽ�*<e��9V�N��TҘ��S\��b&gLB�`V�f�Bɽ�*<e�VJUT�����B���Gk��n*�6%2�c�;�ɽ�*<e�&�Y�"\-��T3�A5�Ǔ:���|��Ar,+�7�Zf�����p����8t������p��O�
�����c���M��l`.��n��X3,Y������ɽ�*<e����
�3O�1�q <�t-*���+.��E��@��ɽ�*<ebMtM��%ֹ�TC�r��b�W]�:����,X�aҥ��A�Y��gu:׈S�y|��5�L/%�
�9�����v��,�����h3�걙�1#Yp�x���]L�EO�
�����c���M�ba�dQW�n��X3,Y�����°��F5�Kȟ4�ЀN�{�?��ɽ�*<eBI�i�ʃ~��0��;�
���"�����n��M����sɽ�*<eWb�"j���5�����N �P����T�O_,���A�Y��gɽ�*<e+�� �{��[��*?}ʊ�C'��u���H�* ɽ�*<eɽ�*<e�[�Aa���=� A6�,붏�#��/9
���ɽ�*<e�L	�^a>��o�["bn
�8CX�aҥ���/9
���ɽ�*<e�E����Ϙɖ����c"bn
�8C	MI{��$�A�Y��gɽ�*<e*��� .5��|y=�M�3pI^C�����p����8t��6nh�
n��8t��}�tؤ�l�k���,(nɽ�*<e��`F�Yt���y�P��8t���ɖY׎�0C���>M"N��b����Rk��.Q3��Ѓ����ڎX8"��ނO`���hA:b=��K�X�[��2�@�pRV���X�E4��,4���?wʉ$�Hl��1�w��A�ɽ�*<e]�H۝��ջ[�ɽ�*<e�, ��T��+(M�e~��V���X����n��r�7�'�\��K��|`	+����p����,��+�k���Q+G��Ts�j������;��"�a�T���`����|C�@D�pRV��x��[���ᦲc�����p�����1�f7���g+ ����,מ
�C'�K��wȖ������,4���?wʉ$�Hl�Y}�c���y�2f!?\��ܰ�AI�/�����n���=#�I����8�)R\�$�}�*U��m<"K����Z����MS������LJ?\��ܰ��|C�@D�pRV���ޡI���+��c����V�uCM?\��ܰ�<D#[hG#��pRV���ޡI���W=CՂ�z�e賙m8E�YZ͆ˎ�kH$E�̽C�6���/��Q3��Ѓ����ڎX8"��ނO�&ѩ�&�Ib��i���sX!�M�����`0�x��\ɽ�*<eI��&6=��a��h���͌:��y8�oh�󫯇ԛ.����cW΀��˺�1�<�Ŵ~T�Y�k���VJUT���Uj+����}NВີ��/�žC���#�N��PH��K�j��.��c�GOR�2��Av�'�B����p���υz4�7-ʣ,Z�'kR�ߴt�D{�	Q}9��݁W/���+�n�/�GAiq��%�f�S��Y4C��uԅs�n �u�HY"���K������n��r�7�'�\ᒺ��A��^��0��N��~�#����ǔ�PH��K�j��.��cۘî����\�r+�=����V�uCM?\��ܰ����_~9����cW����!�����@"G�A�j��.��cۘî���W=CՂ�z�e賙m8E����D�
�RP�8�H���N��P�}r!b&X͸8yw�T�Y�eu�x��*��~�@�"�n�Y��?�0s;��|ޞ<Ĵ�,��.�~�L���m/����!d�<�&MX�a��$\hnA�Y��gmaW�#)�.��QTE�`�/��?���A�Y��gާ������+�f剚l%��K}�����p���ݬ�S��M��ً^����+ƫ��kwO�&뿃BL�\��-���螨c#�jk���,(nɽ�*<e�M��3ֈW��:X1ɽ�*<eL���D�)��b=M�}����微/�žCɽ�*<e��P^}Q���S#��\���V��oޛfe�^C�ɽ�*<eɽ�*<e�{�����u���[m�_xZ��C�ɽ�*<eɽ�*<e���q��Xaa?\��E�h�,�B�r��������-�8wɽ�*<e'$��R��e�����kV�ɽ�*<e��P^}Q���S#��\[-�H���Gޛfe�^C�ɽ�*<eɽ�*<e�!��(�V���.��L��8���qɽ�*<eɽ�*<e���yt�E��G������Y%K.A�Ԋ5OJJ>R}9���}_-.�Ȉ��JrAɽ�*<e��8t������p��ɽ�*<e=@�����W�^a�+���$�K�JПE�[5ɽ�*<eɽ�*<e�*�Ù��:�|��dnZxOm4d�>ɽ�*<eɽ�*<e�)�����w��l�u�ΐdEc�B4�n<6&�ɘ�>R}9���~�9�h��QZ����3��4�����pg���Gɽ�*<eɽ�*<e1��0ɽ�*<e1��0P�7ٝGy�����p���T�t�g��v�'ghI$���.�2֔O�I�_��z�Aj"�3��[$���J�m�Z��~�ݼ-���+���A�2?*�F�s�ɽ�*<e1��d�ߪ�q�7�eC�O�|ˎ���V�uCM+�n�/�G	�y��pWmh��EP$�ɽ�*<e������ ^���=��۩�]5yB=�u�@3/�@�'������p����0ddRy��ҩ�%$����x5��4�b�z�a��Q�:��h�O1>�BɆ��q&�:�e�)f<�a�,x�ń���|s{k�����)Ov,�c���+�f剚��ȇ�}P 쎤d�w�rj9D�m���ҋ\�d�+�ZR�u����Wdꨞ;{Y��
]*ɽ�*<e��;?Q3�0��J����p��AX��'�W��jЭ�w�%LPeBTɽ�*<ef�Æ�=�6�*��Ri�5[�~H���kwO�&뿃BL�\��-����3̧牊I�eC�O�|ˎ�)>˜y/;K���ѡ�p�&h�#�`V�f�Bɽ�*<e`1��w�}���ō�l�Z)^��_������ɽ�*<e�g��-T@��s%��r��\!����ɽ�*<e �)\I��QTE�`�����z0Z/�^5)��ɽ�*<eT��%zؕ��g�q\��/�žCɽ�*<eɚ����堻ۦXI���I���5*�T��W��-���6(xI@�Ŏ� ^���=��۩�]5yB=�u�@3@����^JПE�[5ɽ�*<eɽ�*<e�g��-T@��s%��r���
:��{gɽ�*<eɽ�*<eٞM��EC2;�ZC^��dEc�B4�n<6&�ɘ�>R}9�ܻ�#�ܢBA�Y��gɽ�*<e �)\I�����4����Xo�]�T�s �ɽ�*<eɽ�*<e��<��ݭ�`V�f�Bɽ�*<eɽ�*<e�)�����w�X"��|���@z�Jɽ�*<e'$��R��e�����kV�ɽ�*<e�)�����w�W��-��
�x�*Ӄ�+�f剚l%��K}�����p����8t������p���+�r��y��)�w׽�P�7ٝGy� �.�Qq�*7 ��!J�5!��s7�c,\�|ɽ�*<e�"Uy��\�y!�%��s��LvP���JПE�[5ɽ�*<e�{�����=ڤx*x��^5)��ɽ�*<e����,�4ɽ�*<e����FL�ʻ�ō�j��\�>�z�NSad���5��I�A��;��μ��M��)�Q�o3�� 0n�BA�JПE�[5ɽ�*<e�z�H�?������y�^5)��ɽ�*<e �)\I�����4������չ�<ɽ�*<e �)\I�q����_��P�G"S�NSad����8t���&Nꊓ�Hb�Tw��5�o���6��Ms�������UjA)�q��spoz�X�}��R��Z�J���F�c�q9r�T�?:�;���A��#�P:\����u)�QX^�2���@i"M6f��������5��	"	���?��o��N�1�a�g��ۓyP������1��
O?�p٫j��"�yL�x���Ys�}�q��?Xٵ��5�,����F]�J�������	UQQ*rb�5��6��uF�p�	_�P塙@:/!M_[V�I'�
n� 70^�d�e»�-0^��,�:�	S�uP�M�zK!�g٪�'�)��F�p�	_ى�#�9�$�oWU� ����L�m�C��#��;����B�	?�gwC�N�O�lK���K)��F��P������_#Ǚ��R�����'c.�	?0-� ����Jv���,����@p~�@oH��{T��qɮ����D���,%GJ�=�rW�K�v��|�5������zWG����ʙD�0@]�����>'�6�*�q�t������ϩU�R�4�t������:Wp<!���I��d�>�r=D�9�)�Ί#|�Ӏm��!Q	s>R=��@�wG�ɽ�&���[�O�VG/"���@V��"W���à\j����f���ԝh<K��}|�?�M��\%i�������E�!��o�8���RX<���O��"P)�6�m�`�� P����Y6Z����*y����,��/�&�5K}�*���ՙ��e'�������s�SŠ��z��Qd_No���?�%6=����e���w%fz����I/Ό%��c�q9r�T�?:�;���A��#�P:\����u)�QX^�2���@i�I/Ό%��c�q9���I|�� �V� �s�'�4s�����2s����	k��;l��O����S��mCSfe�%T00�ѐ�ͤ���]����%ޮ+x�(+M%Y�f"h�ۓyP�� m���� Դ��[��Os�w�F��֕pR�Lʉ/[¶���`���c��� �	[�w:���ע��������t��E�̎����D�<L}ڈ�����dn'y&���3��ͨL���K��a9q;���]��e�G<���ߤ#����ө�((|�w��M{� C<�ls���|����䋇�æ��tg������a��4W%��g���$�-�����Mv�'��X�)����qӬ�\ԗ������nx�I��	n�=��ϝ�p:�ɻtpe��IO҅�QҔ�n�zWG����ʙD�0@]�����>'�6�*�q�t������ϩU�R�4�t������:Wp<!���I��d�>�r=D�9�)�Ί#|�Ӏm��!Q	s>R=��@�wG�ɽ�&���[�O�VG/"���@V��"W���à\j����f���ԝh<Kaչ�z�Mf%�l�J�����7N?aJC��B���ڡ��n]h�^�o��p����=����+P
���(�5;B�W��M��v��E�`�w$�P��j�:�mheˣ��:��?Dg,2ms����{Ue#Ty� �I�quȯ����2��ȿ���&�NV����'a�y��2�s�ou_'������`b�j�G���0���-���gpT#o*�L!ˏ�� ֝��*���HCB�7_���7q��QJ�:�����7���<FS����ʢ�� i���[7((�{�!$�w40|2�tF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�dd&1�b���A�3�~(�����\�e^�i�)�9�s��hM�%.v�����u7�~�Mo�gZ�(�*�MK�d��
�B�Ӕ���ս��?Eߕ�?N�$��BU��Gaϯ�J�_��d*��G��[TY�ƪO��{>�E��锠EU��}RfA'����G�3wව�=(�ET`q��Be&�6!�j/xnŅ
F���1�h�ͳu�G��$���_PZ�3�ò�qS��~����!xF2]�J8��tj%��2�-�"���	�c����M��t�-�����^���D٘�S9����7���͞�� $<q��z2���t� ��������]��r9�2"H{�{Vڤ�0�rЯm��a3�S.���*����6k:�S0"槛�`�-�{'��זpx��8T�'N�n�Y.���o�#mL�+}�	�z��E�i�V����U$�k8&GB���;ǩ:]��eQ����s�(�w	���0_PR�4�0$0�/�U��aRh�g�\�hr�ɫ�	��^m���W_�#}y�Cvl�6}Zf���޸��m9��i�S��l��l�VwBG�5�g�)���j��
Y�(t�\"HIV�q�ig��J�}o���O*/��k��$4�
��&�)��^A	�2��۫�FJ���9�e6	̯(HǢ�����h��Gb�f%�e^�i�)�X���*~�2��3vg�8�׮neQ����o]�`oT�z�t��锹��]䯚��gh���D��9��b������ᦼ��� �V���ɽ�*<e7��2B�r ЇA-���$`љR�ɽ�*<e��~^-C�6��2��,`��|��xj.�f��� �3�vo��x���T���j`rc��wo�	h�[��*��`��.��j��e�'T����DSn�*��G;���C���h/����6��I��5�z2���t� ��������]��r9�2"H{�{V��,ǩ6��G�����_=z�Ϯx��p9�,#��*�\���]�~������S%iv��!J�P=3j�ABÓ�z��'}�_��i�RM���������|"ÝW�_����a;���	�P��5����+4G���ȩI%���0Y�P�����\ƴ�u�iޕ "[�*齅B��ǃR�zm�:���sOK�	1��偸����-���+S�D���89~���L��0���:l5��ݦc�AT;��}�C?	���s��D�?R�w�ĝN���hAl3�M�z���+>|�%41�k�a�K~����&�7��cT6�+˿/�!֬9��w�oУ��EE�I��]�@KCս��4�Xn��e'������*�4��f�]���{I�!VʑF�u׊�WE/^��x/�
kEk���f�²[[s=gsO��O�n�p����Q�4�P�X�3��-_�:���ulK���K)��>��]�p�%�e��M��_R5Ƹ����w�xLIo\n�b1$�AZ�jn�-�΢�0�|r�UNp}��J-�4f����/����l�%U�H��ǥQJg�+=�:c*����d��(�ե)f����D���H��n���K�e�~O�=d� ���R��ώO�o��_�^q����y�Gdd`�(�M}�fD�='�w��@/�l�x���Ls�EG,��j��|�#�|d$"���G��(���V���u.`7%<̯:�"fɽ�*<eɽ�*<e��*��ɽ�*<e`j$�v��;'�u��Bb��2[t��	1ÃzBɽ�*<e���!�̿�j������٬+{!$H�K(z=S��Qc�]�<�;B���ÍF��5���5��A�2�W\E|cr/�ӈ�G�3���)��ɽ�*<e�E�"�Z��r��6͡=�W7�mj�O3�O�cZ�ɽ�*<eɽ�*<e��*��ɽ�*<e������G>ܱ�V.S�aB@���:�1���-�O���W����v/zD�H �T?ne�2�K��5���c"��|� -Y3����D�!�����0Y�P��o��N�?�#�4Zc�Ղ�����r�n�Ps�Z��v֨�*@��'��fqr�8���x���Ƒ|ɘ��T[��j0��L�aUX�[\��Ɣ	aLK�Ʇ��՟�Ԕ�p�
���P���Ԭ�ȳ�%-�T���X|xǒ30�ͩ�%��0`��x$��S,؆J��n�fas2
6?��eavg�>�m�L�
0�['ڢA)��D�(q��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8���Ș�v�"�iS{/E�́7�׈�|�.�Q>���ě�T�t�g���i��z�h���}V��|�����N���Q�)y��Ԅ�U@�R#l��=�!��]B|�\��KdiF+N��C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�T�N�:Y�?�>�b�J\�g�gǣJzN+"�s�[L�̛ ݠA�3�~(�Rff��^�:�A����:`�s5n��k�0���ŝ#���0��)�5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8��*���)��Q�k��/ބ�ʉ�-M���*�����K�d��"�_��6�\�u�<T_��5�$�c!��l�)�L��~^-C|��v�&�����)�oXq��hH�]�9i�eE?��]�ֱYZ͆ˎ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)XF#���	��;�?eB*�D��|F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q�ݾ�G�P�!F�����k��TyP}τ���w{�lղ�9�)Y�|6f�aA�X�1�{��F2]�J8�F2]�J8�F2]�J8�~�&T�S���5>�VЪJS5�UC��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�T�N�:Y�?h�!��qF�����k��TyP}�T0�f�|᥀]a���5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�)V ٥�Dk��� V
�,���V�iYZ͆ˎ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)X�yl2���ɽ�*<eɽ�*<e����@��
�ڝ�1�V*h��w��r�!��yl2���ɽ�*<eɽ�*<e�p\�Ì�Q����V����Sk�𷉊����F2]�J8�F2]�J8�F2]�J8�F2]�J8��� �z F7B������RQh��!�X�1�{��F2]�J8�F2]�J8�F2]�J8�~�&T�S��?�Vl��n
��wC��B|�\���CEP�W`c���clS�`M�9�g[����;tF�����k��TyP}�@jk��kŕ�i�S���`KQ���]'E���i
��wC��B|�\���CEP�W`cۓ��:k�UY�s.�|2��rU��F�����k��TyP}�E��C��d�
.��-�����F2]�J8�F2]�J8�F2]�J8�F2]�J8��� �z F7�p��{�$H�4'�{r']n�u�U�i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8��ob���Ow��g�.S��
����c�(g�j&g�jJ���&��/1;7� ����X� �=�;��S��n�P>:�`V�f�Bɽ�*<e�(�[�v��(g�&$QʎÍF��.�f��� ���[`�c���K���P�f�{��t�'$��R��e��䅓�g ������,4���?wS�̦�ːg�K�Bc��v^�%m���� �.?�9��0�[�2AV�f=�[H�o���ɽ�*<e�����Q����clS�H�ס=��0H��r�dZ��8t���ɖY׎��g�H0C���>MX�1�{��F2]�J8�F2]�J8�F2]�J8�~�&T�S��پ� �+�f�LV'>霑�G��rC��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�T�N�:Y�?�Vh��;ko��ܾ����y�b=��K�X�$��-5B����<C����1c���w"�D��O��L]ET�"B|�\�Ȥ`��1�^��z6�V����٤{����p��1I��� !;'�u��B�j�<�9H�?KΕ�qA��V	{�A�W�	 ��lC��We�W��l�S�*�V�'�B�&�Z+����V�uCM�6tH�_��1��=�e賙m8E�04�H����g�H^"f?D����=.{
>�{^E�.苢��w�ɽ�*<e�5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8��l��q�K���)����_�����������#��eۅ��QӚ�E��HgcwX�/����p�������F2]�J8�F2]�J8�F2]�J8�F2]�J8�M��X�{���(�[�v�������7��l�^����.�HX���<��ݭ�`V�f�B�VJUT������F��m��l��s@�ҷb�F���;_!a��܄���d���t�QY#���N�~�*�[g�~�A���`�������Φ����o��A�h�kwO�&뿃M��?�
�1ν�R����)�㪋�k��딟&B��Sh���,��Vx���'m���]�ߔG�=��C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�T�N�:Y�?�h(�(�|8���Z����F�i��J�QMW'�/��	V�v:hc��8D�<kZC��4y��E���0'�����nX�����n��rF2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)XkwO�&뿃M��?�
�@b�?W�5ɽ�*<e($���2��Φ�����0�%��~�*�[gĨ�Q�9 �^,y�J}��ɽ�*<et}ѭN�"��0&��z��n?��� 1߀i��lC��We�0��u�,qS��rT��9���$�Ż.��ݞ�Z��d�
��	D�ܣ{UW,M�d|��5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�)V ٥�Dk�_�4¯c�쨪�I�;s����־�:G�0���B�.��''s\)y�V3n��-Eᩉ�i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8����d��X����G���R�ʹXr�	e���)Cm��Fo�ll�Z)^��_���������M�����ӆ�澮/�žC(`<��"$@����v�S�3���.2P:���[����p���+�r��y��_F��x�J��E|�m;ɽ�*<e��}Gδ�-�xQ��ƛޛfe�^C�ɽ�*<eɽ�*<e�0vsp�x��$���i�S���`p?vT�������ɽ�*<e.�������i�S�����y\@Q���w�*(��Dz�á�X�$���~�*�[g������݊�a^�ɽ�*<eɽ�*<e�ur��!�^�5�E~;�.����֍�q�*|圓��i�S���`KQ��ɽ�*<eɽ�*<e1��0ɽ�*<e��<��ݭ�`V�f�Bɽ�*<e����@��V�T�����^*@�)y�V3n���� ,��I����p��ɽ�*<eO�
�����ƍn�V�+o�����A�ɽ�*<eɽ�*<eU�ʫ�?��4C��n�09W��)!r�J�C��<ښ�2��n�2�)�I�+�'x,�ٻɽ�*<eɽ�*<eɽ�*<e�X�$���~�*�[g#=���U�^yO$�,�ceɽ�*<e'$��R��eU877�P��ɽ�*<eɽ�*<e��5�ex�V���Y�2��a�#���e�3�b<&ygHh�8[Y_�1�B��QT�k�7�M۾����clS��W- x�^�5�E~;�.����֍�NC���&uyɽ�*<eu:׈S�y|��5�L/%ɽ�*<eSE⫄ 2}�-��iD����clS�:�+��[k���,(nɽ�*<eɽ�*<e���clS��W- x�M�J�*�ْ��uɽ�*<eP�7ٝGy�ɽ�*<eP�7ٝGy�ɽ�*<e1��0��H�)v�=E��Rx�5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8���UOZSĥƃ��r`yI`�wb6g�w33@����Қ��Ai�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��8�:o���Vh��;ko��ܾ����y�b=��K�X��M�j�������H��Q�k��/ޕ7~ϓ��;��Ȯlz}��~��WO�"��Ǌ�i�j��'��yl2���+�_���	�?�)ΝM��1����5>˶$1I&��~�af���<(:��?�Vl��n�o���(�2���-}x�9bX�)]�����F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��� �z F7`PP�̥��7���W����~Tʜ[��D���*2-����/�C�� '�]����~S�%�w�V;4�8��	���$�6�l@!	Sv�4��Mk�M�Ju��ќ��ËW^�ɚ�Z\|���o%��OO�X'�в#l���e�b�#�|�9�Rf}Ɩx��NjL�n���YZ͆ˎ� �s���L�b7Tb7n9���S�ڸ��T���'Rɢ����4&��ƞ��f��/ҿ�m�o5���,?��vl-0� �-�R�s��)6�&�z\*�D��|F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q�ݬ4���2�]�"��~p*X".$�����4^�ߨ�G��GB���QX��XW#ƺ�v����?�Vl��n��w��((�H�iˠj&�4�b�z�a�(�[�v��[Ò�����̸���[ �'܄sZ���#h�(�[�v�����L2����`�Q<�@o�L��[��+����+��X�(����~-A�����L$iz'�J_\�ל4�j��h䟒;��������p���j�8]���QOנּә��f���RkR�%eœx���{#OCt-ኂɽ�*<e��^/a�ya ���\ә��f���b&`������VZ�@8r��z�:��
þ6'�� a��4�b�z�a�v��,��T��%zؕ��g�q\$ ��}=K�����p_�ߔG�=��}��Pj���%��Z~��e��W��G�h�
'�(�[�v��-H��5�@��1�_��O�"��Ǌ�^1�5 �3�����,�4����/ַ0���(��A��mt�[�.V`6O|�۾ -`��	�//:����#�>��xl�(T�飳������?ʌ�of�F��i��e��}R�|��W��A��1�����k{��Ty}�zj�"��0��U��j )���.s���2D��%_�y��N�[\��NT��>n.r�P�S��И]h����,��D�se��L���Ӡ��B:l��9q؟��?��6\F�߉�}3z�s"P�A/5���{�)J�ɷ�b���Ւ�tU#�݅�Cs����myW2��KqM�qsdu��&� �r��j%g�*E�Z��(wRET�1�ZAů� ��Ö|�o�l&��H�J�9B�ˎ�U�X���!4��x�ٷ�?��Ŵt� ��R����a��'��FL�j�4F�tˎ3I��(��Hk�p�IwЈ�#oԓ`��Z���GD����4�fgHg)%�RPz
2����$_�>U�V�Q���L�˷P�B�p1����Z��U�`6�!R�4�t���!���8��`�w$�P��j�:�cb�S���mheˣ��|>X,1��>�5T�g�'y{�I��y3AL�����~ָ���}R�|��`iX��-�����I���#^2�}G+�����uP�M�z�ڽS7��v�����
����%�z�M	!��Ɋn�]#�$u�	8'x��)�)�����y�>�t�Jд��߿Kv���������0���L��J���n�+cb�p�f8��H�\=҉7�#�?hX� ]����f�y���WtuZ��ү옊I���R��7�{u���M����飳������?ʌ�of�F��i��e��}R�|��RT�Q��M���W#�(�*� �.6p@�*3d�#_�0!s�,�	���
6�.8�0�T��(�H���-)�|�d!d�H�d�h�ݔ�x��{��õv�̟��������.s����g ��$�L��ow(7ALۗ)��/����0�7��Ǧ��!Fȵa�E�UJ̘�P���W��-�\��\����WgƘc���Jt���M���bf�\c�ꗳ�)�7�;⑤���a,�"�빱x�Q<�^eg��ɂ����c_�o� x/���C $P��!zsv|MC�[��ĺ6
&���?��������Y���i{\�M�Q#�`>�P���=��ϝ�p:�@p~�@oH��{T��qɮ����D���,%GJ�řO���.���C�> f��i��7���x<D� ��U�`6�!R�4�t���!���8��`�w$�P��j�:�cb�S���mheˣ��|>X,1��>�5T�g�'y{�I��y3AL�����~ָ���}R�|��`iX��-�����I���#^2�}G+�����uP�M�z�ڽS7��v�����
����%�z�M	!���=��ϝ�p:�\���YVeX���V�ͤ��075�D����,���AI'�Q�Oﴽ���������
����-��
�=��U&ʀeH��J�	�5!�`G$j`{�+!�Nh�z�{&�@�J˔Qm�4ߟ� �H��K�l�!ڵ?�V�7���Ph���c����:6ݑ��/�׸s7��s�����Ɯ�h�k"(�������j){��	�c/����՝��H\�p�θ��Ɯ�h�Z��g)/x�*B��0�ѡlv���tk���I���v�D�t*�gc�꺉�@jB��Z�!�W�/�Cd�سy�%�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��ې� �r�Z��ٰ��V�A-xE�pxa6oܞ�}h�̠o����Y�u�}�����ˮ��R���E������mF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8���ա8&�o�	rr���6�XoN��5+}4���5�}�'ҺZ�ØK�h%����:�g��7-R��<O7Pג$OJ�7�c��>���DF��t���8����tx�E�Bx�6 �� |���DF��t���x��h�=s���3$A�-���@]�������Y��wAӿ�\pѬl��eZ?��_^�R#l���L�o9Ȃ��_��%l�VV���p~rևv#Z�񋐐��q�撇��SU��~��WT#@�GN�%�mƚ����N&�=�ǚ|6f�aA�����&-�N��)��0]�Ҽ�w	���[�2�R�����d<�s��7Z�yl2�����,#D7��K�am@�nh��@�;��'# &;�J�9��E�M��1����ΦFz]x����Q���.U�[�x�m�������D�U�rfbߘOY�m�� M�C�W��z|���q��<��J%a�<%@p�yl2�����֎��{���\�v�}@'��on~a�2�]ߪF-��7*.E�yl2���Z4�Q*#9O$<�Hˬ� ������;�@��6�J�k#ϸ��F.վ�3��#��'���\Y��پ�?���>��y~JqK����h���b2ޏ�C˾�`,!�� ���J�|�"�����{oۿ/΃�:��c��ѡb� 
��z �W�5��M���E�U-�5"�#F��87U*���gic��ݤ��x��8����		%s��7Z�5��M���E�U-�5� ���	/5��Oh`E�U-�5x����Q���.U�[�x��E�/�k_bLj�]�
�L�`bȇh�!��q!������[<!F �����,��@N7h�!��q�P��Tiy+��VP>�������
v"�+uF-��7*.E�5��M���v��V� j��'�\��}@'��on�fT��I������7-�.U�[�x�3�G��X�5�Ma�-�ORi���D-59N�fY�$����N����R%�16nP|�KU�q�>��1Hc&�>�7�=���EPr�O��aƤû<��q�Iܨ�ֺLl�M��1405C2V�h4W�G�����-3,����n�>n� ��A�׽�Xp�i �;���qRjy�:l�k\H�S���m��E�B[�/.��D�+�q��n�1`s?U�ݱ��g�E�Ի��(R��-�7d{��p���5��F�vc��[��G���N'	V/�Q��6�/�6��gN�梋��N���-��J��3�}ƿMp�Z�������
v"�+u�@b�%�S<��1���F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��KM��b_�~G7@��H�2':d����H�NLa��b`��S�`TJ�+t*&�x$w��,*�+��ă�d�K^�T�*k�Sŋ-���V��bnz��d�vu4�o�i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��1���`s��jxg�����l
nb��g��X��S�q����j}/��}?��.�w <>k�Z�<�]ɘ]�0����r���3=�x	c(��H������3��N�]��I��y���]N���3���J�0�v���3">/eJR�k�/eJR�k�/eJR�k�/eJR�k�/eJR�k�/eJR�k�/eJR�k���S)�uш��t�d������#��������9������m[1^m/eJR�k�/eJR�k�/eJR�k�/eJR�k�/eJR�k�/eJR�k�/eJR�k�s��4�}����p����Aך��{FI�-tCa��R�ĖhԷ~��0�mZ �/eJR�k�/eJR�k�/eJR�k�/eJR�k�/eJR�k�/eJR�k��U{]%�U)e�YJ�h�W 7(x��"��,A�!#JI@�V<\[2>�sA��/eJR�k�/eJR�k�/eJR�k�/eJR�k�/eJR�k�/eJR�k�/eJR�k��MN�)7L'uQ }\�e���0��E'6a�����D/���/�j3:�F/eJR�k�/eJR�k�/eJR�k�/eJR�k�/eJR�k�/eJR�k�/eJR�k�1y��1wjVA�Y��g;��n�l�D�E���M���'��x�	��������2/eJR�k�/eJR�k�/eJR�k�/eJR�k�/eJR�k�/eJR�k�"M�VyQ�K�P��m�ʚU$`v�Zp&�Fr�>����)/�zC�~��T7��S�/eJR�k�/eJR�k�/eJR�k�/eJR�k�/eJR�k�/eJR�k��U{]%�/�g���ɽ�*<e��Ň�;�$l
nb��g��X��S�q���.D����Lf��/eJR�k�/eJR�k�/eJR�k�/eJR�k�/eJR�k�/eJR�k���I�,�Z@�NSad��D4��*6�v�I��y���]N���3���J�0�v���3">/eJR�k�/eJR�k�/eJR�k�/eJR�k�/eJR�k�/eJR�k�1y��1wjVɘ#�7���ш��t�d��@��	ʔ�������9������m[1^m/eJR�k�/eJR�k�/eJR�k�/eJR�k�/eJR�k�/eJR�k�"M�VyQ���(�r������p���k�\�!�g�>����m�X��S�q���.D����Lf��/eJR�k�/eJR�k�/eJR�k�/eJR�k�/eJR�k�/eJR�k�/eJR�k̵��Sv�7�U�e���В�S����	�Dh��n�Ad.[��S��J�Ub)�'��b
��w�0�z���^A+�o�$3��4��e��:�A`��Cr�mD�����K~u�p̍�>��L�&�-���3�]3pkx��LV��і>�F��d��`�bJ�Ub)�'*8M�`��S?�1e@��^�(�Ѳ1�8���gADpz�X�	��Q"�I�g��{�t�X�%%�KC�qo������5)�>ʻ��5c}?�F�#�5`��)���}5�K#�7;RML�}y���2M� b5,�Im7�@�����8	���)��P*(�1񷊑�o�I�G��Q���F;���!�)I ��������W<Q򒥩��}��`���Yr���W��ʤ��&�u�ƾ�Ź����޵	�p�3W�����g{G�Pxף$��:g�`�M�>3��h���!�O���ʄ���tn�~٬3� �$�f�J������$Ym��� u$�%���P��:S��]��Q{��%��))Z"�he$���뗊:�g��7-E�U�ֻ405C2V�)�s*UB� <Е�_6��[@B�=9����r���̗�	Q�������Z�&dH
,�-��j��h���<Q1�������Y�c�9Ձ׌�:Ycq��6^��J�q��_0�e�0��S��xߕ*�v�=<�x�u�O�:><JGc�cG�$��;��SK�54��`԰kS��<���S�2�w��8��	�D�_d�Ǹ���Mb?ߎ��#��M\�[�#\|/�@�^M�yWeS:S��]��[a'��EqdRn_�_�z���s�O���8	����e�o���=LU[$"��م�S]��ʣ�G�Ge�;)�m�9��H�ty�A��?#��#Ia�.GD�dz�Q�Ƨ���:��2k������!���K�<Y��^~V����/���?�䵓L6 ��\�e5�:��T� }�t�\#����r��>|>�^�j����-��P��
�,�d6���y���d�n:`_q�>��1H|�r�����A����f� n�T����-��G����2��W$�fUsWW ��Gt�$� f���_��l��Qc���a�
:�<-�:NF{��V̴�c䙵1c�ȹ[�0��S��P���5o��yvyr���O��9��\
����u���y�ҝ[��R�lȏg�����L<ިgA�+�����a���o\h��4mS��R��b���,�|U��0}�6�,H��ݺ�� )�hk���k 3�'�)���.$�k� �����L�	�׃2��!�(I�8��U�ٰ���˫�l�������#���@$v2 ����w�� R2Y[v�_��7���~y�x:j��QbZ]�Վ3� 鰫@ވO� ���vTX���}`K�	�;޺�v�*ҹw^� /ϭ���~���b���7�r\��%[P�=<Fz�5�5�Ma�-�O�)*�Qy������03'�u���A��աD�,d�\�&�cK��� �Gseݯ^k���I起ҝK
'>~
Z��A>��'P^�й��w�s��8�?1/<��sш-�:NF{���Y>��ۂ�}grj���5�F��B)d�[k�ƀE��m�ΐ�s�m�	hT{�[�$vY$P9T��4�p��&�;!��)�c�Ԛ�/��=��I��ٰ���˫�D�l6��)ԋ�N#(�/��>4��}bV�3�@uzwZ������)��6��O�s�&�;!��Zĩ�O���Z��^�*څ��}�t�7��lEXФ6��4t��lݮй	s>R=��@�=K8no��u �W_DפT��pVCø��A�Z��k���R�I]�!Unt3hT�)����NV<}�OhI��� 1��o��u��5��j�A�0���d2�3�(�J#��X���W#R��p�uC�E!͠aX��y�5꿨��]̙[���-VԬQ"���{�Fw����L�zHm^�,OD�aUyP��9`%���VJi� xN��zf�7۬&�Oe�v;�I_4\��=-$Bf��46��+���X��0]����
O__	ꅱ3"�_��+�-���1׶0W�X��c���{�W{l�0�H;�c�>�q�	�`�����B�2`>�P����p��S	��-�:NF{��7��<����|��vǿ)���)�e��v��L�p�	�WO4��rg�U��o�:g�p��Bpq[I ���Hv@�%�C_�SƤml�ǀ)NY�ھ�I��g	2�3�m����"?��Р���N��i�˘ڇ
�܎[��s�Ի�	>���ey t[Wn�.�/;�Ua�.GD�dz���A�-+_cj�c�Y[v�_� �7��r�uF@��Gb������a�Ɯ#�<��׈H+4�������NxL �?&ħ�3�O�/��KbY[v�_��N!
�bl^#z�R�au��;�=�h�b\�(���7NZ����r/����˕Gjp�|�н@�1~���C�)�-�:NF{������T��21�f �xB�� �7��r���W#QR���<E�/�����|�:�#�Z\#ہA#�R�t^$O&��XXv�-�	ª�ѝ�U(a�jy�yQBX�k{sAa#�pnZ.��k�a[���y���6��)ʯ��~��f��\*���m��Z4�Q*#9�t���Y[ԯ�	�c/����՝���;�O��	W/�b Ar��{v���Δ��B����W/�p.�q��	�c/����՝���;�O��83��K�����ovL>��\[����q�0���_�Tk���s��#V�,������u�#l�g�hre;_��f>4yR/�������q�0���U�^�(}!�LڜY1���.�d��p�����Hh�P�?N�M�#ȲsU�n���0x�)�x��mM�mʘ�F�,O�H�ՖI����Ӵml�ǀ)NQ���X�4oCƞ�Xܳ=ܵm�_��?��{�h?���r��c����hQspB�-�r������0x�)�x��mM�mʘ�F�,O�~J||Q֟z���4��92U?c���:�����)�1l�Vk�'r-�N�~)�X��*����n4C<!!�DIB�� ������߃D���u<@B�LY��1{�:���]�*;�@��6�JCȸ7�}�d��p�����Hhߨ�o����ŗ��]+��q�Qy[�^Nђx� Ή�+��c������+�(�T	����YT�������l҆��c�]~��P|c /�ъ��HRe���1H�����q�>��1H���s��r�[�֥Z��!+��}�w	��Q�~\#����r�"7'汦|�o�	y�p�?���7#��80���h&� ͞����E�Ի��(���NY����A�a�jL������Q�E�8#��@��v���iğ��!q���Ę�S��PG��t�8��Z�b�P�g�0N'u�n��}�ebEв�E�u�+��P�����~`��r���#p%b�)ʯ��~�vŬ!	�:Nw��Ҩ7�T�4ˁ��}3����k�����d����p��=F9��V�N��<�")C�Ѝ��7]T��{�!��}3�����3�N8��T���s8���.
�_F��D��k��-�)>˜y/;�)%��b0��a/v�sݏ#P�Q�K�\UcjoAh�q�`V�f�B ^���F�d��p�����Hh�^�(��I_��NSad��wL =���R����������L�8j�!Yn��R�P�7ٝGy��_F��x�J��E|�m;����@��R͞��V��a��{e��S��]&^�H�m?�G�NX�Jj�*^�45R��K��/�žC7� ؗ����Pj�Ʌ'5&7.�٥2���o+z�������8�^����? ��9;��H��}.A�+g�ۉ���!����M��,B8�A���
���c}n��{lL���գ�����	�����P�g�0N'u�n��}�ebE�2��4���A�Y��g�P�g�0N'u�n�O�{<i~3�ƾ��e湷^�6C_ZWA�Y��gf�{��t�ɽ�*<e���g�q\��/�žC��
����@\�y4�R���5"&���Q��`V�f�Bɽ�*<e�Q}g��ml�ǀ)NQ���X�4oCƞ�Xܳ�p#����d��p�����Hhߨ�o����(r�ǝ_`w4:p��ɽ�*<e�	�F��ml�ǀ)NQ���X�4oCƞ�Xܳ��{Ŵ`t�}3������E~L@ɽ�*<e�/���%�C�Ѝ��7]��Ǩ�������KN�䉲����ɽ�*<e�+�r��y�ɽ�*<e���g�q\TD��;1��f
�#O�������,z�w.@�|������ $�Y�gɽ�*<ewL =���R����������L�8j�W�B|^�(��s�ԧ(}��ӧ��4f�6i�ɽ�*<e����n��r'���7�<#�o��-kEMއ)d"�����FR8��?K�6�`��R��\Y��پ�?|��5�L/%�VJUT���\��M��O�*6x�ˈCVE�OjN���0x�)�x��mM�m-��:�"���
:��{gɽ�*<e�+�r��y�u:׈S�y|��5�L/%�+�r��y�����,�4��7S��N5�*N�s!������4Nvc�����X��:�g��7-�9�a��d�"j�
]55�*N�s!������>֠د�	�c/����՝�����
���2����� ���������MXD��$NZnx�ԩ�����U�{u������с����^	>A?�wT�X�\��3�#<O��
D�s����CU��S�#��;���U͝�N.���Y ����	�X��x�N.���Y ��-���.nw2�V0�w��N.���Y �'�=�3��J�n��V�~�c�9h�W/�p.�qi��3�)�*���s�g�����)iyz�# �X>F�UA|�܇���`���D{h!嵯� G���M`��l�4�k-���F(\��S&������uu�M�#�¡��'�K����B�z6�#��Ut(�.O�� !;�g�^T��ׯ��l�M��1d��dZ}eR���N[3�Y��e�����YT�80���h&� ؝����@��Mˡ늙���t�kB��g(���JU�p��{�����P�:2]�$B� HsEA�#q\Z����9�l�h������c�^-��`e!�J�ߢΨ�Lv���S�?(o�c^���,�fZ3)��L���Ԉ�  5˃"�Ѱ=��|����480���h&� ؝����7��N�tX�$�(?R0�ڊ[߇�Z,���3�����
�tT�0^�5f����eQ���j�h��Hk���}V��yzXƻ�2��gƧ)����y4z����X��x�N.���Y �C3���c{[-:�x6� d9���n'�����kV��!��(�VcZ�c��d"�^ϭU:d��KaH �5ɽ�*<e��^/a�"ڀ#�e�P�F���jX�'�>Q�b;!�����N��)��pN.���Y ��NNeͩ ɽ�*<e�epG5�xP�)qOm�~�c�9h��d�5t4��u�û�236�C(4}g=s���3$M�7�'~ɽ�*<e��^/a�"ڀ#�e�P�F���jX�'�>Q�b;�P��Ti9�:�9KU�����{T_���F��aE�gP�djJu���e�gܓ�f�{��t��_F��x�J��E|�m;ɽ�*<e��^/a�"ڀ#�e�P�F���jX�'�>Q�b;�P��Ti�	�NV�^F�Um�����u�û�2�X
�ɰ�f�{��t�����/ַƭ7X>��'4M���//�%
q�sڝ�o� }�uKO��m2T ��c%�`V�f�B��}Gδ�-��$Q����x���]L�E�Q}g��ml�ǀ)NY�ھ�I�m}S+g�/�~)��B���^�%����1bdY�Do�
�0�C�y-�l]E? ��9;�q���\u��\�r+�=�ޛfe�^C��CVE�OjN���0x�)�x��mM�m6�U6q{�A
ߔD��<���������d4�1�K=�y�Ԯ{T_��ÅU�c���$}[)<P�7ٝGy��v��,���(�[�v��[��zz^5�|835� gsӣ�j
a��vM���'��x��l����o:%���j�&��K��5�@ kK�׋He4r�dQ�h�͝�����Q��/��7�J&K6������&q��`n������d`�50izoO� ��5~M���ӏ��,��ːKU[���'{�b�Ӗ�)$��x=ëjs��_h􆗟��+W�L��W�X�u.im�o���)ʯ��~�08O{F+��[������d|��a�H��E�y-�l]E? ��9;ȓ�K���֨2+k�ݓ��n��`� ^���F�d��p�n��5�u�o��\.Ȥ�tQ��]D�$NZnx�ԩ����e��b l~Rp��4z�{�����F��j�Bʨ.��t���B�bl�acuiE��7ۅ���z�%̗��w���\͠�l������R���`�a�4Cf�g��΀�Do��P�/��2pؒml�ǀ)NY�ھ�IؑS�P�5 +�0����epX�q�����/J�!#�]0;�G�	�M��)�atBҷ��c A�[f�矑��ӆ�澮/�žCݕGء����a/v�sݏ����p����	�c/����՝�����
���2�� ;@���!Yn��R�P�7ٝGy��_F��x�J��E|�m;����@��R͞��VTO�Ɩ�tz�S��]&^���Z�|�[JПE�[5�CVE�OjN���0x�)�x��mM�m6�U6q{&�vg+)��m�>5��U0N'u�n�Q�>����Jۿ�ғ��G���p���b�!�!����M�UDF6u�r��O�u�W����I|�k���,(n����n��rwL =���R���`�a�4Cf�g��΀��������,4���?w�+O�[5��b����2������3�	�}վ6��]��ɐ$]0s �>fRĂ�m��ɽ�*<ek�m�&.ǖɽ�*<eU3�=�dJПE�[5�VJUT��șC_�SƤml�ǀ)NY�ھ�IؑS�P�5 +ݳR����Nɽ�*<e7��{�����	�c/����՝�����
���2�� ;@�ⱕ���3�	�}վ6��]��ɐ$]0s �>fRĂ�m��ɽ�*<ek�m�&.ǖu:׈S�y1bdY�Db�Tw���*�wC`�}����*X�ZF�i���l��MM�X��s��弨���'���7�`�M�ެ�z* Fp�2�S���7��׽�hq���T)�}�xۜ��Fs(iɗI"����+l�	ܛ�8P��VEmm'�]ӟ�0�����-nU��Gi
��Cj����,��@�h'r��Ay�A��/��po���=?kV��='v���c>9��Q}g��ml�ǀ)NY�ھ�I�m}S+g�/��m�˗�g�ml�ǀ)NY�ھ�IؑS�P�5 +�/�)#�Gi
��Cj�R�W��3N�܇���`��X���)���L� l%n[q�Qy[�^Nђx� Ή��g�E	�$�3����~a�2�]ߪ�q��
�6����\�UF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�HE��޻'�j�/>wH�éa�G/�8?���N�k����r���Ǐr�b1�Z��	#;e�p�25�Ǔ��N��߆�B�bQ�]��1Iثhe�k�}8���kƶP.yt��xl�	<W�N�&����L���5����OR����j��o\#����r���W�~�վN�p�����R��AS��<���!��T�:�_%aG"�,6Z���9�=�z���b��-{�HFrE3qͿ5���f�7���1��~ =�f��&ak9�o�F׼�C^*�6�m�K�am@�~��M��r��O�u⇪	[Wd"�rt(��o�d���|��+��pb5}߽C�M��-�<�������Q�����^EG5�td'QZv�i��`MlZp
T�m�B����GjP; X0N'u�n��}�ebE���d4;r~Z�K���0��f�M�
V8��+ Z;��N+ށ|M��t+c��T�=!�KE�8#��@��v���iq�Qy[�^N�!7���V���g���>y	J�X쟋�^tD���ÙEǛ'�=�����������u�#l�g�hry��$W��(���6;Ѽ���d�D-{����%/�����M�����`	���f}��S��i�nP|�KU���^G6A�×,3a[�ZG�N�6鯷���B;W��o� ӥ�bg6��W�q�>��1H��
��	�~(���`�/eV�W�P��o܆��eo��HI����{s}��{��T�.h�+��յ˄5�p��iZ��t�	��%O1�'I"lt0w�C=[�ђx� Ή���m&�� ̠o����A��K��hp��Ԁ�F�Y���~N���C�.sK�s(�?A�Ҏ&�Ё?m�-�,�X�Ÿ�f�2_B@�~%.DI���:��t�%2�/	J��hא�܇*9�2�\c�5��u|R���GX��a��Xڟ3�8�H�d�h���� I���}�t�wI'[]
*�J���oE����:��C�$k5p!,�7ڐ9� ��h��'i沃�Z}����Hc�9�%�\T|Aů� �B�#��t�(a�����z}�E!Ͽ���!Lؒ&�bL�.��. ����lB��,zyj���0_��A�\��B�N��%졖*��j)?��(a�����@��$�G#�ӵI�0��#Ҟ�s�-I@>������BP�\_�0'���I"ʈ�W�rB�������i0aXK��2��H����D���i�6 ��Z�)a��\ `L���c��}W�R�#C,��n�Yx���|��/_��P��r�k���g��� H]K�s��K���{T��
�7`�	�6�#'	��m�:��eH��J�	��[W�DC�"�N�?�ot�'��#~D��\��KB����VL��'�s���7K�f*���b�0qK�s��D�1d�	!4wI�o P��z9����D�����e�mu���H��H�
:��p��؋9i�^��,1DԾ����\J���H�.'a:�s�c�A �Ы���VI#�1z���x�q��Ǝ�b\[��½�#��$̆���5��0^v�'-�r�D��6�^i~��b!�t�&��9W����z��\(uՍ�N9T�k���ՏZ=��7�^��j�4ִ��2�������W����j){��:eLE7)�پ������8B`}��?�(��G���0��L
�(��7DJq f�&�'F���Ϫ0��!�4B�7_���7���2�fo�����7��?��L@��m:�(4�����[7((�����6�IYt���$͛Jm�X���F2]�J8�F2]�J8�F2]�J8�F2]�J8��ې���X ���5�<����������V�zBB��Mg��S�+��hcу����Nk_���D2��j��\�ra޵D!*m��HK��5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�4)�}Uh����n�r�Z�}=��8��z�S�M:1A�Pɔ=Y3����j){��:eLE7)�پ������8B`}�wG��L�qC��ଡ଼�F2]�J8�F2]�J8�.��A�5Ȟ�|���	����й���*�D��|F2]�J8�F2]�J8��5�� �ۍc���<	�4,2�
Y[Òfɽ�*<er���4GH_�.ťw� 9�]�:�H�T��qɽ�*<e�^6bD�k�/{���lӎiC��WH���ɽ�*<e �2p0,�����O�4�S�?ߐ��&zl��z;� v��S�iy�눽�A�O@";\��� �sDDL	��D2��Wu|Pr���<�&f�u�_�$�!��y��s�r���4GH`I���=�*e����D�fVA�0 yɽ�*<e}aՑ���g�H�Z�g� 3傈Moɽ�*<er���4GH�y��d��J�_�p!%?F�ɽ�*<e��Ec]���ڤw�_�T����h�C �G?�L��r���4GHJu�e��릟:K�i��t���J}E�ɽ�*<ex+����~����S�Z�:���B�p�?�r���4GHS�S�����tgv
�i�S�DJɽ�*<e�`�?y?�<���y憾~�c�9hfVA�0 yr���4GH�a&+.���cr�j�����k�:?o
ɽ�*<eV8��	�D�<���y憒E�I6�L	��D2r���4GH�q=�J��P�"�YZ/�ԂA�ɽ�*<em�ZG��v���<�&f��MS�����ɽ�*<er���4GH�ɴ^����øxQ@Q�;H�T��qɽ�*<eg�W�g��q<���y�.�w <>k��h4���r���4GH.��rى+cr�j���5k:e�."ɽ�*<eCA6eR=�<���y�
鿤ｮ�h4���r���4GH`aٛ+npcr�j���Q�6>q�ɽ�*<eQQm�:��Mڤw�_�T�
��d��	B�v5���E�r���4GHd_� �	�\�`�P�J��wP��9�ɽ�*<e4��� �
ڤw�_�T�"�#$W&��L�0Ō^ܛk�$-���:��\�`�P�J�����G��Zɽ�*<eą��bs�ڤw�_�T�o���R�-�	F��ݏ�r���4GHU��r�\�`�P�J�ܒ��5H�ɽ�*<eJ���=� �!	�{�`�RR`jɽ�*<er���4GH�⌨�g|@6�����H�T��qɽ�*<e.<]�8{Nb(X(i��5r����9!ɽ�*<e�߄��a3�k�/{���m����kH�T��qɽ�*<e�V�w��~e�>��9�B��K�ɽ�*<e���*[���8g��$���F�+Sxɽ�*<er���4GH��{}.`�� �P1s�j݇�M�uɽ�*<e{*o��^�%1�M�@���á���ɽ�*<eh�� пAț���DsN��8H��!���pXb�sb�[��,*k3Ӷo�`n�L�T'r��Q8��;�#��l�
�mal���{}.�\	�je�1���b2ޏ� �G?�L���paË;��o�ˆ����<l]j^a[���K��r���4GHO��.��h���*b���]iLɽ�*<e0�Bn�gNs@�'���>R}9�ܲ��]iLɽ�*<e�d8E��,�����F2]�J8�~�&T�S�)�o��Ymo��E�"�DEuyf��C��ଡ଼�F2]�J8�F2]�J8������Q�onv>�v2DaZqOW��_��_�{���S��ɽ�*<eɽ�*<e���������En�]H��Q1����Dh�GW����Q�q'{�ჭ�u�l�֐M#zlp������5�C"R�R��!��DEiɽ�*<es]�� ��%�W��)��N� �7oJ�o�Hnτ�����&2}��$sN��8H��r���4GHK|�t�9u$���$t�_rw���+h�� пC}�/��cF2]�J8�F2]�J8�&���y����JY�?�4h�� �DZ�	�:����8�5����fF2]�J8�$�䠢O)X����9|-�ჭ�u�lo���@�I��� ����~�ڹV���ި}E](�N���['@�(-�]�x�����y�>3!��9��Δ��B���t��R(C�%���Nbq��D��Aț���D��~�1�7���,��!	�bđ;z��dI c:��iTS�Z�:���?K��qAț���D/Χ��,z�r���4GH�USm��]�t��R(C���j���3K�['@�(��3�Գڸtx�E�Bx3!��9�؎��홓��h_��'��1=?ض�cAț���D��~sEr���4GH-�]�x�f�5~��r:9y����?K��qAț���DE׭#��
�r���4GHe�>��9�1$$8d v9��A��ݩ2�('�Aț���D�$(�d¼��@��p�q���@	��p�q�1��ŧ�ۥ�{}.���:^��x�,������fk�|B�����b2ޏ�t��R(C��J��}�e�;�$�D�^�<{������F2]�J8�~�&T�S�۵����0��m��yQ����Ci�ܛ�|�F2]�J8�	C7��3�^��� ��#*ɽ�*<eɽ�*<e:j���+�0�]�{�;�5����_k`ɽ�*<eɽ�*<e��_��l�.�+:-nP�5����fF2]�J8�$�䠢O)Xe�����%�U�q%PKԭ���zi�ễ��X�1�{��F2]�J8�����q�ݭQc���øxQ@Q�;T�F-�U3^MͿ���q���
���2H�ڸ��P��B�a�h�ɽ�*<eɽ�*<e��9�Y�X�o�D�m�U�\�I;���ɽ�*<eɽ�*<eMͿ���q�r���-��~��W��XgM�] �YJ�D`�����)-:E�q����d��yN�F�8I����N���*��H4.��_M���5@��*kaMy�P����g�d�8�72L%hQQ��p��u��dɽ�*<e{��<Ia���rq��&(�xt��:[�Kn�:Ou
����.ɽ�*<eMͿ���q��P�6;7}q�cW����yl2���
�P������7k��/��:��$���-rvT-�Ǆ�@확yl2����e��i�Y����L�N��T�F-�U3^�lև4[@.Qu2T!�ҕyl2���ɽ�*<eɽ�*<eɽ�*<e���$;�����K�,���a->�d�wo�	h�[ɽ�*<eɽ�*<e�u��=���-��P������9��,��H�!g�ɽ�*<e:�]�,VD��v�i}�"�Zr%��������a3mɽ�*<eɽ�*<e��;@�M6L{���V��'x�|���C}�/��cF2]�J8�F2]�J8�&���y�����:_���@�bY���l�VUQ�F2]�J8�F2]�J8��"嘶�������9��ɽ�*<eɽ�*<eĳ���|w�ac]8���}����N���Ϯ���O�)��A���&@��w@��4�(y�5��M�����x��{ɽ�*<eɽ�*<eB��1_�m�B���	��y��:.H.�4&ꬶ�Rɽ�*<e´T�&H�Z���<���^:{��ſ5����_k`ɽ�*<eɽ�*<eL��M?��q����6��9*�D��|F2]�J8�F2]�J8������MP���A��<3�X�b]ъ����F2]�J8�~�&T�S��yl2���ɽ�*<eɽ�*<eɽ�*<em�x�˝��zxʯ�ؾe��|)��A����:��$�V>�Vȅ�J�_����z A��hAU6]?���i�m`�+M֏��_��K�`H�ڸ��P��B�a�h�ɽ�*<eɽ�*<e��3��>}��!�(I�=LU[$"\�I;���ɽ�*<eɽ�*<e�ub����"vЅ\�P�TT�I����N���6����=�ɽ�*<evS+ё@���ɃH�)S�Y��*i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)X�'yP9�������V��C��N��-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��KVة����C>��M �IꜦ�4�ݝ���&�|�D����H`.A7�+i�����K	t�nQ�ɽ�*<eOM1���s�"B��l�-׍d���fo)�J<��Cq�g�k	,�{s~��Mھi��͗
G�H\�ߢP��A;�����l���zA�Y��g	/�`*\M}�˃Ng��q���u:׈S�y�է '����ۓyP��vߦaJ��V�E7J,Zݪ+i%��f�V�2=��ǬH�[����=HI~����`n��i� ]���ow�����O����s�c��������W|�B�6eL�v�k��S�1�V���z���.4W�jՇ���5��b��\Qi<S����㢒mԳ=c@�LTP�@+�1�7 -����sEK��]�3�־�b��Z�4�?�k��S�1�V���z��.�w <>k���� 
���H���N�Xw���[��~[CLO��/e��u�x�&C��L`���Θ��mCߦ�o� :����*��q%'cX�K�X����z��B���"K��w�It�Ke�%zQ�P�W3~K�R��N����t{2ۀHj\��k��vR�K+^(�s��s��5���
�N̝ V������C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�&���y���u9~8)f.��Ռ��gP�׬JCR��H�.�т5�K|f�mCI�^�Z�X��*�ʪl�VUQ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^PXq��l����T0�q�(�[�v����ioK�C<v'�k�,�Ntk�3<ìKV?��˾�[(S����㢒mԳ����с8�ie���f������S��گI�V���P��Ti����o�����с8�ie������ϊɽ�*<er���4GHe���+�I݌U��]�¾��:^����bQ�ƮP�]�磐$�S��=�)��L>���b2ޏ���F�<��O�;8W�fT�F-�U3^'�=�3���lza���הܰ&���R�5�z�%�F�}$[f ȿ�0������X̽�ި}E](�.�����ݤ���{.���xXi+}�S�axVX�1�{��F2]�J8�F2]�J8�F2]�J8�~�&T�S��勉:=Ȑ���9�J�_�w�'T\��?�n�z�# �X>�$N��Ϯz�q�f�Lw�Z�l	������a��cp��a?�le�I,H��ݺ��	CǑ����0F�d=;h�-���*�D��|F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q�݌U��]��:���Y�w�u��V|���8����O��>M�K�ŷ���".$���Ę�c� ��Y�ϤM���m{��v].����p��}��Pj�	[QI��)pg~z�|g��w��'�ɽ�*<e1V��3m���4��j)�0�V-�~ы�VFY��d�{�s&�N�d�>���%qX�8Zl(A�Y��g1��0�����n�x���]L�E(��Î�HXM궿?(6�U6q{W�@iO4��޹f�^@Dp �q�cd{�T��%z�:�[��P�X��X���l�VUQ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^�b�ё�R�Ï,h��P�.��jI~�z��`um=�4�i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8��s8���s%����3JПE�[5�>6�`G���b��M&ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eލ�6���iԙ�&�Vb-���Ծ����.ޛ�ih�~��ɽ�*<eɽ�*<eɽ�*<eW���W�~ ɕ?kV7��CÁ�� ��B	�D�������L���tgv
�G���c�]��G��8��ɽ�*<eɽ�*<eX���b��)_��D ��b2;�*�e���s%fd��<�]a����l��B	�D�������L���tgv
�G���c�]�?����ɽ�*<eɽ�*<e&� !;��"CGͭ/��ɽ�*<e����n��r���n�U���F\�U�ӭۿ�d�a�C�e|X���F�<���4�d���h4�:��cD�~�c�9huFS��4�r���4GH�{T_���!Bx��i��7'r��ѫ��P��Ti�	�NV�����s�g�4�1��
�H�8�H�c��h4�:��cD�E�I6�'*F�l����*���lև4[@n�k���Yiԙ�&�Vb-���Ծ�6�_� �n� :�t�[s#y&cɽ�*<eɽ�*<eW���W�~ 6�U6q{y���P���B	�D�������L\�`�P�J�vl��%I��bR ��Yɽ�*<eɽ�*<e&� !;��"_xZ��C��g�4�1��וۏ�`ǌ�����S�Ƃ��ɽ�*<eɽ�*<e��*����W-�AzA�Y��g>�m!Y�
��
���t�U�Y "�t��{d�.{KP�^�%ɽ�*<eYS�\*_���ċ�d��?�k��p���b�!��e|X�0��W�d��`�_q���ɽ�*<eɽ�*<eɽ�*<er���4GH���|�ʃ��B	�D�������L\�`�P�J��`-��}!ɽ�*<eɽ�*<eɽ�*<e��R��Wٷ ��㼽|liԙ�&�Vb-���Ծ��#��V�;0c���]:ɽ�*<eɽ�*<eɽ�*<eW���W�~ �V�A���&�R������=��Zw<Tl��0�g�4�1��{�u�~O{��r&�F6�����'*F�l��ɽ�*<e��*��Y�=�5G�������L��M?��qpx�����m����k��݄�L������Nj�S�Ƃ��ɽ�*<e	��LM?���W��#T���޶(:�e|X���F�<��O�;8W�f��݄�L�������Q���>m\0c�r���4GH�J&K6�^Q��4��xL��M?��qpx������JFV-O�;8W�f��݄�L��)*z�8$h�#��IJ<��PI������/H�(��K���P��e|X���F�<��8r��c���݄�L��5��77��	����r���4GH���"�����=��B	�D�������Lv9��A���1��';U�����L��uFS��4�ɽ�*<e�i�ɱ�*ey0�z �}Hk�K{�ԵT�F-�U3^A�Y��g>�m!Y�+�r<5�5H�n�?Y':��w6�ݗ��0�:
�'*F�l�����g)Y+��NSad���e|X��#�z���&�-�WK*e����D�uFS��4�ɽ�*<er���4GH�<�6��R�im�i�>N����s�g�4�1������İ��K���1�����ɤɽ�*<eɽ�*<e��*����z�Z�nG��.s�x_
��`�+VMr2����u�_�$�!�ќ�+nR]���h����%��������jw[�x./�j��>6�`G�t�ؠ0v3>�Fv|�dU�Ӥ"G���d$s�:B�S�?ߐA�b��0��ލ�6���MͿ���q��P�6;7}49�iv (ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�#ȯ\�N�px����Z�-��K#d$s�:B�ؠ�ʔ*O�
����KvB�"��A���=��Z޴h�>8�?�ER�WV)ڬ�����{ɽ�*<e����m�Է���2�������LtV��^���>�A*����?t)̶tV��^���>�A*��B�.�ǧ�o�_F��x�gƧ)����ך^!NH7N3�����,�s�]�{{�v��,��*�D��|F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q�ݯ��`�?�
�t%Է�dz9��yy\X�1�{��F2]�J8�F2]�J8�F2]�J8�~�&T�S��E�40��dYAzN�!�u�"J�z�6|"��K�;��μ��M��)����n��d��)%��b0��a/v�sݏ��Ę�c�����N�ھi��͗
�`�"5F���rq��&�caT,ҝ/0H��r�dZAN$(��5ɽ�*<e�ڧ�N)&���9���.�>Ƒ�������
����ɽB�kj`▘9�E����_H2x���]L�E�8{����hT^)�����ߔG�=��ɀ����[:Vjӧj�lrj��`�^��ӕS�q��J}�Ĺg>��fU��ɽ�*<e[-?F�^��\���
�9����k2�G�CzU��e���K�9�9��`V�f�B��|ޞ<�6�M���:��C�n�����h3��.
�_F��D��k��-O��V�n�&T ��c%�`V�f�Bɽ�*<eݕGء����a/v�sݏ����p���´�'V�5�e� �zy.2P:���[����p������,�4'$��R��e��䅓�g ����� �
�������,a��ߗ� �P�� j�Z��JПE�[5ɽ�*<e�´�'V�5�e� �zyM�3pI^C�����p��ɽ�*<e��cw�<B���<���^��c��d6ɽ�*<e�J�@1�췆�Z8��H
E#LPA�Y��gu:׈S�y|��5�L/%f�{��t���8t���ߔG�=��h��]L�ދF��ݕٰ���˫�4i��
U�a�e��^/a��I��,i�K�am@�n�M���r����c`yX��_�Ԟ�Y'��˾�[(#��z�Z�4�?��SCR'3����Z\�J��E|�m;*3ZC�q���^����"�#F��8�⠡�����-�8w�j�8]���'������<���^�V7��ɳ�f�1��e�+�r��y�Q���'�}�ٔ^qt��5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8������MP��J��3��)�?�B��_d�Ǹ���Mb?ߎ��5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8���n�.:�	~���`V�f�B�z�a�{�sSu���eɽ�*<e9{�z�0rMͿ���q��P�6;7}�~�p[�3�Ӆ��E�N*3ZC�q�f@��S�c��.�$� �a�=Շ�A�Y��gZQ�R�"=:�1���-��ڧ�N)&���9��k�h7T�������Y��
���61^�L�֎%;���͢^\w�i��k,�
��
���
EÎe?j¸�`�T�ɽ�*<eY�=�5G��f�y��HZ$��Nnpm�x�˝����`�7.\�zu�V����kwO�&뿃y�P����g����!�p��u։�ɿHd����ߔG�=��n�������~�T�ȭL>m���8�ba�X-�.[G����p�����]��q�-���Ծ�{`is3Z�em({�):��m����kfZsh��g�����p��{��<Ia��/���?��f�2N�2���NSad���+�r��y���H�)v�=E��Rx�06vk�&�ީ�q�Go?�CmM_M���D"��
D��H���/T� ���\����q�:�P��#�p4�`���J���F�c�q9���I|�� �V� �s�'�4s�����2s����	k��;l��O����S��mCSfe�%T00�ѐ�ͤ���]����%ޮ+x�(+M%Y�f"h�ۓyP�� m���� Դ��[��Os�w��*CM�.S���bc+Ji �8s����6e���%���2"��
��4N;L�Oc]����m���x�?���wIF��E��OU���2ޔ��e�����{�n�q�r/<��\�D?('h(�m�W�K.j\�NIf���'Q+j���p�D;&��'��K�����c�׈�}���	'��@Ybs����Q����N�?�9�LZu��,�K���G.|DT����(PЎ��=H��|�j�Y�ٰ����DlWIo)��87��ݥ&�@O-�
pΟ�����Ȼ��*���ՙ��˂����ɪ��H����I��	n�7�q�BH�������(�k�T���cD�HM��נ#s��3��.5�)(�/��>4�S{v^�F��MF�R�i�LP%o/LA�\��B�1U�<`<�a[��6����J��N͝�E�Z4��������7N?>����R�����z#9m
���������h�>K	�K�7	�j����m%p7m�R���|"ÝW�qe�
��Q ǂ�L5��k���g+��jj�h��#B3�q�2�w{8����y��Z��Vof�*�D���K0Sj�����ޑⳮ3f�d
��v�g˨�&�;���`j�{=�}\��8B`}��?�(��G���0��L
�(�D��}L�,4��l�ג$OJ�7�
�`L�=�CeL�f�ZSl�Ȅ�{ڪ0��!�41ҕ�G�9����DC�#�/e�x�P�f��H�H�i�YEK�x7^LX�1�{��F2]�J8�F2]�J8�F2]�J8�~�&T�S�?%6g?��q����ޓtd�X�$�H+�ɚ
��
>o�r^�������P��_N��^��v])�rta���D9$õ�@�Z'�8z�L�Y�l���c��J��&�+{${K}Ԧ
�W�ʤL��ً�X;_ړ���C������phl%��A�
<�>��r�&;1ɇz(E�I�;��FCv�w>�5� ����13+!D>� uA�6[��G���;��b#�x��\��9�(���=�p_(PX^1�[~%��A�
$��rL�F2]�J8�F2]�J8�F2]�J8�F2]�J8�
�c���z��g:�Bح������A	s���B�p��3Ԅ���.�?g_[X��S �����
l�Ma��͙]�ͻlU�� <�ZBgM,�Q�.#�5��jnΨ�\E9;�J�+��V��0��E���ޘ ~��fɽ�*<e��*���l����m:~���J�^*���ɽ�*<e��*���l�����'Z�Qln�5Ǔ��G�tx�E�Bx��*��eZ?��_^��e���>sK�EbcW����]iLr���4GH��j|�$WM�|]:؄��ޘ ~��fɽ�*<er���4GH	�&���b�P#���n�5Ǔ��G�tx�E�Bxr���4GH�؇���Gk����n��r8�K���VĤ�n���_N]y�<z���;�X�8��*�LX�ɽ�*<e�M+DW��l V{��������׳2�����(i��;k.nHw^�����<pb�L�׏�����ATV�6J����*�������%�4�-�I�M$-����Bɽ�*<er���4GH7�C�!#% mOu�r}��aO�!�ɽ�*<e̧th���ĕ��cW�&2}��$R�����aO�!�F�O�e�wW6Н��d=MK(�b�ɽ�*<eɽ�*<e���*[����7)Y�8O���>Sp�ޞx�-�ɽ�*<e�a�s�f�N]y�<z�\�j׸'��^Hɽ�*<e{*o��^l V{�����g���.�Dz�.�ɽ�*<eHw^��肳�n2q���ô���M�|C�f���� x��FF�[�[֙Ζ4R���*|3k.sb}Hi�X&�M��aO�!� ��J�e7ڨM!Q��yu")�
B�dC�r��ɽ�*<e{*o��^⃦�q����D����Y]�9"���c��Nz�wج[�:Gc/���Θy�i���_Q��'�nL�n삾=Y���rh���=�d�~p��z�!r_Q��'�nL�n삾=Y����F�i<]7�C�!#% a����_Zf3�����S��ɟ����~^-C���cW��Gk/�(�@�c�`��bT�>�@�3��)i/��Y��{T�_0���ɽ�*<eɽ�*<eɽ�*<e�l��m	�yl2���RKD�vQFɽ�*<eɽ�*<eɽ�*<e��^O�f�x5�;M�����ב��6%J� �<�?x����f����N���6����=�ɽ�*<eɽ�*<e�6���	Nb�F���<ȑZr%��������a3mɽ�*<eɽ�*<eɽ�*<er~�F��[��eh{q������9�օ=�v'���ޘ ~��fw�u��V|�����~.O�~�e�U�5��M���(�_W�k�6ڸ�OB���c��LL�cw�u��V|�W��J.Qu2T!�қ5��M����W�����Dt���/B���5���w�u��V|�(.%�,�Ǆ�@홛5��M����W�����D�uۨ�T~�;�K���S�Ƃ���ܚ����&P�_������W<:KRKD�vQFɽ�*<eɽ�*<e���F+lB�#����Zr%������S���)�ɽ�*<eɽ�*<eɽ�*<e��u�%�㗟��<�E��
�a��{T�_0���ɽ�*<eɽ�*<eɽ�*<en�$Ӝ�>@���:܎��X��]�LN\=�)��#�Ε�@g��*Kv�6���	Ny�P����g�p��U�p(W'4�l&ꬶ�Rɽ�*<eɽ�*<e!�4@�+/���?��=��c��v��~��W����Zɽ�*<eɽ�*<e���F+ZQ�R�"=�S��O�yl2���E+��I���:��$ɽ�*<eɽ�*<e,{�&ZԨqCƧ.��X��]��zN�����ɽ�*<eɽ�*<e�6���	Nf@��S�c��.�$� %`���;��e�����%�U�q%P��N��#��̻U��Xp�$�28 �f�[>���ɽ�*<eɽ�*<eɽ�*<e��9�Y�X�o�D�m�U�]�9i�eE�p��u��dɽ�*<eɽ�*<e{��<Ia�������X��]�LN\=�)��yu")�
B�~�;�K��>a��b�����
���2H�ڸ��P���S���)�!���dT�4V{1�E��D���Ȫ}�0)�||�,�h{�a->�d�W�����Dڸ�OB���c��LL�cw�u��V|�lև4[@.Qu2T!�ҕyl2�������=н��5V���E��D�ɽ�*<eq����d��yN�F�8I�X��]��zN�����ɽ�*<eɽ�*<eMͿ���q��/�]� FY:(|��1�yl2���RKD�vQFɽ�*<eɽ�*<eɽ�*<e����UO`TeE+�O✜�\-�F=��~��W����Zɽ�*<eɽ�*<ekwO�&뿃,�M����yl2���RKD�vQFɽ�*<eɽ�*<eɽ�*<ec®p"�.bt�2"���~��W����Zɽ�*<eɽ�*<ekwO�&뿃���t�i��Ͱ�1��׿��~��W����Zɽ�*<eɽ�*<ekwO�&뿃K`m�B��<�� �[i{T�_0�����a�;^<0H���i�z��Y��`�11�}J�5�vӸ=].���W<:KRKD�vQFɽ�*<eɽ�*<ekwO�&뿃y�P����g�.�?:.�f�Zr%��������a3mɽ�*<eɽ�*<eɽ�*<eLݴ��;'�u��B�Zr%������l�*�g��*Kvɽ�*<eɽ�*<e����m��qCƧ.�����N���6����=�ɽ�*<eɽ�*<eMͿ���qp)2���@�h2uvm���7ޮ=c@�LTP�@+�1#�s%��5�'�q�Z�-G"v:���x�F�ud�^�~���㿷�JYw�8�r�rz���~N�|�9ݱcI"	@��IgL��X"/�$�Q����Ì����V��+Er��f�<Q����Ì_Zf3����n�$h�����~2�"�&��y�2 �9bA��7�����?Zݪ+i��dd^�jb�~3?7`�n�n������F��ע�]�nO��~3?7`�Z�=^�ć�~N�|�9ݱcI"e��%��п���P�7�ow���X
�Q�onv>�v�j��_�6=[ALt�^I���;�X�\�rd5�ݖ�9��^���9��!tQ�onv>�v�3��0k��S�1����Sf�e'%��@�|7��s�ƨ��h�v�BЈ�Q�7�K:6;E��V�B�ލÇ2a?zF�`�v�*\ɹ��~i��&���ow��?�c�y% �9bA����;�X�ͨeD��qڸ�OB���c��LL�c�X��f�漯���l�Hi�X&�Mo�H!�|�G�S�#���C�L��-<��pN�3h�2�A&&"�hA� ˯nkB�JݗX��?�`Ȁ��?jx�.��k���-@<�/���x\��斳q4I�\6���ҥ���Qw; ^ӭ+Ј�Q�7�s-�1r��?��OsN�cnNMG����P���74���{�@@x\��斳��H�J�Tx���L�N���]]��.��=HI~��:<_�U����vMk�~ы�V �9bA����;�X侮�Z���{nr�����p�A�������UJK����pZe'%��@�|���ɗdW�Ј�Q�7�c�Z��U!@Qj/��<N�8���\�yu")�
B�#�3֟Ӕ ˯nkB�J����=f��ҥ���Q@�đ�k��S�#��k�]0��A*�fJ����)-��s�m]��ȋ�D�Y�_���=HI~><8{��gk�]0��A�o_�|\���onJn�5Ǔ��G���P(���=HI~����`n��k�]0��A�o_�|\�=r��֯��"��+�~��ԧ$���i�'�2�5��Oh`������<���;��oX��Ę�c��J��y�Ih.!%��*
���|H�Pk���,(n�����I��UD��S$ɽ�*<e���5p�bF���|��р�������A�Y��gwp���	JПE�[5ɽ�*<e��M]!#5�S�-qdy�@Oל�:�L����`��Q������v�M=�ɽ�*<eq)�_�������Z��ɽ�*<e�+�r��y�f�{��t��9߿GE��>�I��t|{�U�K-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�T�N�:Y�?S��6��
�3w�E�?����#��(ՠ��Xի���1���/<��Ђ]���b�Q�p4�8��m?*�b	Z�2v"�eSTI~T�إ��Kˉ�)�)W�gmr�YZ͆ˎ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q������2�f3�I�z�c�����p���D8=�m�4�!���A�Y��gQ���֧.o�\�1��/nɽ�*<eJПE�[5ɽ�*<e��ٛ�ɣ�����p��I�[��Y��AR4=�������p����-6L#�T�I+v�y~����1⾮/�žCɽ�*<e㕬�ph���%W��	q�ho?ɽ�*<e�z���^B~C���#؟K�]�ɽ�*<eP�7ٝGy�ɽ�*<e1��0��S����	DX~[�=�ۓyP����I*㏘�(���	��F��7 Z�عK��!�W��\Z)�4�p���b�!��`V�f�Bɽ�*<ee���3�IA�Y��g�/�o��줣�dM-��9�؆�p���b�!כ+�r��y���S����	o���p�{��=�u��5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q���t�R����H�E���s&n�:|1�j�1����(Jʰ^��)��@�j�M�(�bJR�4�c��U��l!�!��Ҧ �l�C���,B�:��1�Z��'(�^��q�ѽX
wپ��eE1���i�uX̑�OO�X'�Ͷ>�8QV�������^=����D�(�0@��{�\��?�n�z�# �X>R�+lDb��	==e�PI���?�G�׉ .|����`L&���7)�
ǃ�X���W�P��R�+lDb�n�a�c�EG�ś�ӸM�PP(P�Gb)��W�g���%�#VCHr�~�%e�FG�V��"d�����2F�e��ʵ[�B���ZD�c
.�4R�nZ< #M��X����8Ni�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~E�L�JC��_�����%��0��P�줆�׻;��O�t�� Y䏏NAI|3k.sb}Hi�X&�MMj��*2j�n�5Ǔ��GD�>�V:!���QĥW����с޻���
n�5Ǔ��GD�>�V:�q8���kAF����>.����`�E�	ah����ó�$��L�X���=HI~�'cǬE�|�M@��j/��I����u
����.ɽ�*<eɽ�*<e�&�|�D���Ȅ���g<u��rnN�-����4ud��E�p��u��dɽ�*<eɽ�*<e� 7maH��mA��4��&[�ߌ鼮��~B��<}Ex ˯nkB�J-�̮�F5��'`���C���8����5I	&�5�*N�s��}�ʳk����V��+�E��D�?1���A��˾�[(����ҥяL�8H���bd�e�
*�I:�h�w�W6(C.�����- �*���m������1H��z$�Ķ�l�VUQ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�.��߮p���~�|�Ԛ���t���-��F!R�0t����dY�!�*�D��|F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S��(�[�v��Ls!�EŬB�$DW���W�~ i���!�)��p��r��U���f����Д�٪,#�=^XOV�3yn�3��Q�\9R}��Pj籐�^#�DhY��F�����"T+h�����Æխ��A��S���Γ1��#�s�#�3w@�㗟��<�Eq�Qy[�^N�<�h5�\��T-��|�YS�\*_�m��F�e;_��f>cHZ��r�8;7v������$�\o=��O����ö�#5F��2Y�"ey�P����g����!���O9�))���z�IYLy��+�`ڊ����F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^}Vo1�(��x�9�b�y�_�܎��5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q��(���|�b��^�i���������fuh�+�fKˍʔ��j��ej���/iԣ�֎%;����\FGMͿ���q������4(�R n��ŕI�(^��(�nf�:�]�,VDژڇ
�܎[��O9�))�T���N�LZ��Ę�c�H�h����\�()�Ľ�6�6�Ok���,(n{��<Ia�����(�-����)P�hxf�}��Fʪp)2���@�h2uv<�WV
v��Y�tѥE��䅓�g ��������9�Y�X�Nl�>*�2�G���_D�y��ej���8t��0.d�չ�R�l�VUQ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��瓂�a!ca���ɔd����u!{W7f'�:G�/�ݠ�zY��mnr*�p��S	���)�<A"X�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��Mh���Wn���tQ<[����您�6���	N��HN�E�*�V+��9������"`#�V#eν~�/�lޠ�
���T��Ӯ�C�����N�IC��fH߷���F+���8������"�yu")�
B���tA�������萑ںy�#�)f)-�m8րJ7�}�$�:�x�9yu")�
B���tA�������萑ںy�#�)f)-�m�w�E}�tؤ�l�k���,(n%ߒ#@Nܱ��
���2e�Hu/���ҥ���Q�C�QS{Ԃf'6qGZ i���Q@Qj/��<N>���#n.�������z��#�W����.�yu")�
B�K�]=��"م�v��G3����s����,�4���Ɔ��"�����F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^����D�����$��� ��;��vPm���C��7��� A}�l�VUQ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��s8���s%����3JПE�[5!�4@�+�[�eonD	��/�Gj��E�	ah����ó�b��cJ�%�ט#�i7J8�Kj��m쩔R[�%��iՑ%�hP���.9�W���m�ˎ�%`x���]L�E�6���	N���,(Q'�Y_f��_ 楁2�s�m]��ȋ�e�#.�'H�sN��
����i˔�[Ԉ���L�N��w���[��~����p��%ߒ#@Nܫ�D�\å��`��^��\N4HQ*�fJ���ߚ�%����ٺW��X)�5�*`��h�(�3J)�H��rgz�i9�����\N4HQ*�fJ���ߚ�%����ٺW��X)�5�*`���r��s��
A�Y��gwp���	JПE�[5ɽ�*<e?1���A��˾�[(����ѿ�!��;�X謁�2�]ʳ�$�8B�h8�y�#M^��P��D�\å�1
�T�w���L�N��������b/Q�onv>�v�5��rj7��XPWG�-*�5fx'$��R��e�����kV��+�r��y�9�ݞR��=�5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q��x*ّ�9 �`�cr�vB.r�7@B��d�r'� �>=w:��5���0)�m�9�L�#�W�E<\G�-�j�he���+!٢�`3q�7�¬뤴��%���P�� $���C��n.wg��=�SD<�l�VUQ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��v�����UV�ː�	�*\ɹ��@��*kaM���l��y����K!�����с޻���
n�5Ǔ��G-�̮�F55n�Q}6hA�X����}�n���5�*N�s��}�ʳk����V��+P�]�磐$��˾�[(�EX<�"�I� Ů��*����n4C���ӕ�6A�X���~Y��a7xL�#�W�E<t1���U��:��[�[�W+S$��n�5Ǔ��G-�̮�F5H ܷD�҄(���|�b��^�i�������L\�� D�>�Li�D���HN�E�zo��.�%ߒ#@Nܫ�D�\å4�и5֪]���,(Q'�Y_f��_�4�b�z�a�L��̽.�,\Pش��M{a����x�^6��u���S���,\Pش��M{a����x�^6��n���`;��7�������#m���n�h� 	�`V�f�Bɽ�*<eL\�� D���b��V�o��O��}�n���ɽ�*<e�#;����w_�}�X"n�^żH�P��`��m٤ ��S�o���8t��0.d�չ�R�v����0��[{���F��ױ0�N���~�o ��ghfB)v��V"�4�y�0QV ˯nkB�J-�̮�F5gV�3&�����?�'��pG�3������с�=�v'���ޘ ~��fw�u��V|� ����(��^Xj�?�����D�
2��C0M`��l�ݯ�b��B���Zx�c��|�M{ ���d]7�q/���	��b׎� "�k���,(nO�
�����xV�����k@y�<}�F�~3�?~e'%��@�|F����ޛfe�^C�ɽ�*<e��^/a�|�2�GL���?�'�8h�u[�K,T��pj6�U6q{�3��NW�yu")�
B���py��Je�O� ��C��z(��CyO ˯nkB�J�W/�p.�qyO$�,�cekwO�&뿃%�-�b�fwC�O��ƀQmmT³�p��S	�ȟEX<�"�I���Z~���� �,�P"~(<���s>�o����3�=h�`	lq74M!d�>����g4�L����p������,�4'$��R��e��䅓�g ������(��Î�HX��M�d2��F�a_�-r]�fe+O��ż?�3����HN�E���?%6�Ј�Q�7驁/�r���9�J�a�D�~3?7`���M|=�GL\�� D�{&eRW|��~N�|�9ݱcI"�J�XlE�x�(ZZ,^F��O�R5�+ұ��{-�-_���Umj�A���Hyk�Ck���+h���dyO$�,�cekwO�&뿃%�-�b�fwC�O��ƀQmmT³�p��S	�ȟEX<�"�I���Z~����ޘ ~��fV�H�*K�Aؖ��!������Ȗ�q:��sTd�1Ҋ��&�r�FT:�^�P.q`�5F���&͂8ik��w�|����N*-�7�L���
EФ�2F�y]�Xd]7�q&3x��kNe)��J_����;<ɽ�*<e�+�r��y�f�{��t��_F��x�J��E|�m;ɽ�*<e�����Q�v�]l @$W��4Րl^a�=������8���V��v	��Je�O� ��C��z(��CyO ˯nkB�JD�>�V:��e�gܓ�(��Î�HX��M�d2�ߙ�8�{E�K7�H��o��O����~�),��Je�O� ��C��z(��CyO ˯nkB�JD�>�V:��e�gܓ�f�{��t�����/ַƭ7X>��'4M���//�%
q�s��Kv�V��P1޸���$Q����x���]L�E3ƹq�nNs�]�|tֿk���,(n��
����V�݀��Ε�\��I,�s�]�{{ ^���F۴�˾�[(�EX<�"�I !U���*./�j�T��%zؕ��g�q\��/�žC�cǭ�����1Ҋ��&�s�B�9� 6�U6q{����r�A�Y��g�~�x���A�X�����DQ���v��Rc���J�EL�cm��aOr0c�/T��-���ߔG�=��$ÞXu5ȼ�ݝ{w�� 3��;x�J�u�CK�❕y�L��Y@��A��ghfB���j;�����p��O�
����d�l9���Eg2������`V�f�Bɽ�*<eL�r��NB�o��O�;UT���2ԃhL�ە�pfy������޶(:ɽ�*<e'5�_�����`��m٤�ڨk�n3ꇝC��&Q�onv>�v�u@�@�ҝ�:�h�W��J�J�b�l�I{d�!Y�ɽ�*<e��<��ݭ�`V�f�Bɽ�*<eL�r��NB�o��O�;UT���2�{V�B�n>�8jdH��^Xj�?��ɽ�*<e�CVE�OjNJ�EL�cm��aOr0c������c�!��J�EL�cm+�;+	��"�_엘������_�A�Y��gu:׈S�y|��5�L/%�Y�tѥEo�
�0�C����YuI��/�]� � uV�-8�������3w*����`V�f�Bɽ�*<e���ð1�jZQ�R�"=�&�AD��JПE�[5ɽ�*<e��
����V�݀��Ε�\��I���Kj���pG�3������p��ɽ�*<e�[�eonD]8�>b=��ŗ��]+��~�n�k9)����g9G�C�.�B&�#K�qj�	`�<���!��v��j��ɽ�*<e1��0��8t���&Nꊓ�Hb�Tw���Au���T�]0;�G�	�M��)����n��d��)%��b0��a/v�sݏ��Ę�c�����N�ޛfe�^C�ɽ�*<e�߀h[j����y�\�I]8�9��Ψ�\!����CVE�OjN��y�\�I]8�9��Ψ�\!����T��%zؕ��g�q\��/�žC��}Gδ�-���YuI�A������s �� fW�ܹ �Ivc��u��L�[�`cl��lN����� �
�������=9 <�t-*�ޛfe�^C�ɽ�*<eO@����vc��u��L�[�`�:����\�rɳ'ԙɽ�*<e��<��ݭ�`V�f�Bɽ�*<eC!m�C��L��Y@��A��ghfB���Q6V��NSad��'$��R��e�����kV�T��%z�s����+�1���:(d�a��	)/�zC�~��_/갛�~s�L9=ޛfe�^C�ɽ�*<e��}Gδ�-Ek�ꬊ�Eg2������`V�f�Bɽ�*<e ^���F۲F���H�.zat���y�Pɽ�*<e�q�И�mJ��E|�m;ɽ�*<e�CVE�OjN��y�\�I]8�9��Ψ��
:��{gɽ�*<e����,�4'$��R��e�����kV��+�r��y�9�ݞR��=�5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q����fR}]GZ)]�u��&�j�d���MD��GrX�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��Mh���Wn�]0;�G�	�M��)����n��d��)%��b0��a/v�sݏ��Ę�c�����N�ھi��͗
ۓ]d�����j3��a{E�6��h#A�Y��g���g�q\��/�žC��ky�-��g�`C���ƥ,`��u������r�s�C#e�uO�
����0�]�[��B#�<	ݽ�L{���"ɽ�*<e����1H�]�ڽ1
s'0E�ft� <�t-*�h)VM��''��2\���l��`��M�L>�;>clϚ�y�f�NSad�� �.�Qq�*{8[v걡���r1K]dz��%�'"5�7d��_d�Ǹ��״��w��/۔�	�H�{֧`�]�h\@{ޅ{�c۔/�C�t �ţd�6�#�Eɽ�*<e�]qJ:��ď��\�JqM�3pI^C��&Nꊓ�H��Gm�X���N��cJ�A��!�(�g�`C��̔A��*��k2�G�Cz��5Vq$��ô���M�|C�f���� x��F��$^��*3ZC�q�"�9u��夣�P1޸�l�Ik�yl�m��Fo�ll�Z)^��_������3ƹq�nNsd�p�{nɽ�*<e��`V�;�.�j3��a{E�6��h#A�Y��gwp���	JПE�[5ɽ�*<e��`V�;�.�j3��ac�ٮ:���ɽ�*<eEk�ꬊ�(H��u�6�9c�lC������p��%ߒ#@N�Ǉ�P"�!J�I \��9�����J�M��B迸Ψ������>���AtZQ@uk�T'$��R��e�����kV��+�r��y��+4YZxx�X��X���s8���s%����3JПE�[5Y_���7M�L>�;>c�	* �����R���76��&.�;sO�
����]��]��7��I�tsC��R}%�AD��`V�f�Bɽ�*<eZQ�R�"=:�1���-�r~�F��[�Ndb��`n�D�P"������%e�܉���k�i���R���7��}�;��P�7ٝGy���Ę�cxL��.��gry�,�ߺ�0����Ű��x���]L�EMͿ���q��R���7=�����ɽ�*<em��GB��'��2\�ȃ�m��'O�_d�Ǹ���M��9ɽ�*<e�-�YR����- ��m�I���7����C�Ȩ_�b���S����R���7���@A0,f��?4�ď��\�Jq�B迸Ψ�mb��Z�1��rɳ'ԙ�
�9����O�
����b��4ڠ8��UC
��W�e�e�:x���]L�EMͿ���q��R���7����}&�EA�Y��g3��֪��(���9�ri�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�&���y���JG�?�>���#8W{%�Kn�:Oy��RÂ�n�>��	)�S�ee��U�7�A1��d�7�Z<e�6~JV5	�Á�Cߠ�L>,�:����L��()`u�R}c�X�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��Mh���Wn���tQ<[����您�6���	N�]kKE���=М����\!����!�4@�+] �4r�\�f�	���_xZ��C��U�y�$�"�l��Z=؃�	���A�Y��gfMT�Ҁ��0�,c ʣ�M6ʄRRg��Ę�cR;P�5��N��I-����Lz�������%�hP���Q��q��`V�f�Bɽ�*<em��GB��'��2\��|U����'Ĺ�`�7.\�P�7ٝGy��)�w׽�����@��H�h���N~�;N��k���,(nɽ�*<e�ܚ���ԃi*jZ�+q����d�A�Y��gf�{��t���8t��}�tؤ�l�k���,(nO�
����.�N&��w᠃ж��Q��q��`V�f�Bɽ�*<e�-�YR����- �e��L�
��Mh�]=^j���w��O�F��:ɽ�*<er~�F��[˨|L��N1���|�ʃ�����p��r�֏��9��H��cx&2}��$�r:_ʴ��,��V#x���]L�Eɽ�*<e�?T ]^�;Ѯ�Y�=�5G��޶(:���F+T kq��B�۵���n�
��nE��$�<��sٔS 4X����p��r�֏��9�1A���-�q��q�"ώ�ߊG�Yua�N~�;N��k���,(nɽ�*<e�ܚ���ԃi*jZ�+q����d�A�Y��g�6���	N�bd�e�
*:�L|j� ies�g�w�:'$��R��e�����kV����Ɔ��"��}Gδ�-&2}��$R���8\h2�5ɽ�*<er~�F��[�,���gXS�4z�d��%��d0�b�1�g�`C��̹�`�7.\�zu�V���জ�F+��)�<�;��O9�))�e:M��H���Ę�cxL��.��gry�,�ߺ�0���˽훖�ʌ&�]���%ߒ#@Nܥ�&��tEd�?T ]�����6���ŕI�(^��(�nf�!�4@�+b
��*)D�ܚ���ԎMK�g��,f��?4ɴ{�'�c� 0.d�չ�R�l�VUQ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�]oE���n@Q����_~`"��1׮�w�'T*�D��|F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S����(E��:�ũb�\�G�9������/J�!#���tQ<[����您��
������G��a���_���\=��/�žC�̃n	���7����C�Ȩ_�ai^�73������g����HU��T��8t��}�tؤ�l�k���,(n� 7maH��mA��4��&[�ߌ鼂�q�Q���ܚ���Կ��)�5��Y�G����'3��.&[�ߌ鼮��~B�f�{��t��
�9����'4M���//�%
q�sڝ�o� }�uKO��m2T ��c%�`V�f�BO�
�����GbY�%�JПE�[5'$��R��e�ũb�\�G�9���{E�6��h#A�Y��g��<��ݭ�`V�f�Bɽ�*<e�� ����7����C�Ȩ_����=:v�P����9�OM�L>�;>cy��6�ɽ�*<e���2cm�Ӗc��<���N:�r�C
�V[� �.�Qq�*�izO�j��R���7���2�|ɽ�*<e�#b����>&[�ߌ�@5��c筌ũb�\�G�9���A�Y��gAN$(��5ɽ�*<eZGjr�7+����g���N��S%���@z�J��8t��0.d�չ�R�l�VUQ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�]oE���n@<u��rnN�-��S1�WT�C�D֚LR�5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q��1���|[ ���%[J<Z�F�Aܘ�t�� �?�N lB
~� t2	���!;�'d����e��d�Ej��A)�^U�[��a.�Sl܍�P���QRM�I2'�=�3��Z������U���al!�d�`�I�)i@)��6:3�h|�;Z�ހl+����Z���#�������7�g
�hV��GAv&0%�F�1����`"�Q��#Y�܃M�*����n4CT:�e�����U���alQ6z4£�ӑu������,(Q'�Y_f��_�lo�')�(z���`���4Ӗ5}��Pj[��a.�Sl܍�P���QRM�I2��F�=�����g9G�C�.�B&�\�K�����kN:>�_�!�V��������Q�����-�L��װ�|�B��eTq�����M���r�	��d�p�6 }my�V�O��ML%)��},��Ul/�U�Y����d���;��O+�Ó�Q;ge�{�ƙ�v��~��Q�YC��/�žCpK�FB��F�$��]!�#lѥ��_���\=��/�žC�̃n	���7�������#m��)/�zC�~�9��b����#m��^Ń���\��&Nꊓ�HL�"۠��JПE�[5����@���ݝ{w�� 3��;x�J�u�CKxP�:���X$m2����YuI��/�]� ��;`Ǉj��G���d�a��	)/�zC�~d]C6K�X��� 3��;x�J�u�CK���j}����,�4���Ɔ��"�"Uy��\�V�W�v#@CH5x�`{ѕ5��l)Ȟ 胨RJПE�[5��}Gδ�-��$Q����x���]L�Eu:׈S�y ���%[J<Z�F�Aܘ��'1QC\��\!����T��%zؕ��g�q\��/�žCZGjr�7+�� 3��;x�J�u�CK8�[S�7e ���%[J<Z�F�Aܘ�t�� �?�N����@��js���J�U���al��ٸ.1Y�v��	�A�Ղ��9���y��{��R��/�+;k���,(nɽ�*<e���2cm��d�p�6 }m��ī|���^5)��ɽ�*<e�+�r��y��ŕI�(^$�7¹Z7�q����d�)f���7����C�Ȩ_�+b�:�#a�������u:׈S�y ���%[J<Z�F�Aܘ��'1QC\���
:��{g'$��R��e�����kV��+�r��y�9�ݞR��=x�N����!*�,;E��O��]�Q_.e5i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�HE��޻'�6�&�9�X�����=��>[�$�Ǐѹ����Z�R|���^�ҝ[��R�ɽ�*<e������T걥;��E��=��>[+#����1�Q���=����M2uƐڙ���;����Í�:�ԃ��2�j¶���D����ˬ�r����/��5$�c#z4�����,��JC�Ȩ_��L����Ѷ���#m����tχQ�Y[v�_�ɽ�*<efCc�!���p�ܔ"I��Nb9;�3-�Q�6q=$'�R�	6҆ی���2~b�>6�X������sT��~ M�4��ṥ �uv���h���"(����_���,%1%���ښ����h���NM{9q��ؕ+�qz?9]R]���%�W�����ByZ�������^�
:T�{��*UWY��ÁM��۠�VP,5ya0C���B�4���;m*=ֿӏ�
j�34?
���Z6F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8���e�̣Lݴ�����ȉ=��4ud��E߄ǲ�:	S�9�%�^�}De�<����W-�Az;��OG*��[�[]�&8�0��4ɕ?kV7��vM��������jЈ�Q�7�^MXm�VU�	(�� ���l��y*���m������]v��sK�EbcW��F��P��`������J�8'p^x�#5�*N�sڸ�OB��|�E3�̟@���[�eonD<��s(꺒��9�%2��_M���5���?�M���9�Y�X��ڄ�}n�lv�dF4��"�9u��夣�P1޸��tf�� r']_�@[��]�|tֿk���,(n���M�����ӆ�澮/�žCY_���7M�L>�;>c��!G���vE{��l�./�j�kwO�&뿃M4U�|?�iP��[Pɽ�*<e��B�������p���11�}J�4�-1,&'tɽ�*<es��l�sȯ��L���{��<Ia�����Z�Rɽ�*<eɽ�*<e�!Yn��R�ɽ�*<ec®p"�.R_-�5M?ɽ�*<e`�P?��A�Y��g* ����2,�IM�+�I����WU��x��F!,�s�]�{{MͿ���q���
���23�&z	���ɽ�*<e���tU��ɽ�*<e���-rvT-��P��'ɽ�*<ef���{�+��NSad������2J�EL�cm6D�ά/{vE{��l�./�j�kwO�&뿃�l�06���Ҧs��xɽ�*<e��B����&Nꊓ�HL�"۠��JПE�[5kwO�&뿃�jHi���7�+���ɽ�*<e�:����N��rq��&�k0���MͿ���q�8ߜ�R�ɽ�*<eɽ�*<e�B�LJFU/͛���0�kwO�&뿃�wH��[�ɽ�*<eɽ�*<e�:����Nes�g�w�:kwO�&뿃%6m�gɽ�*<eɽ�*<e�:����N�~�;5��kwO�&뿃��0ך�������\�wɽ�*<e�:����N�_�av"�5�1�ذ{��<Ia��ɕ?kV7�#奯h�ŗɽ�*<e���W�o,�IM�+�IF�������VU�	(�� ���l��yɽ�*<evE{��l�޹f�^@Dp �q�cd{�kwO�&뿃������J��Y[�9Aɽ�*<e�:����N���g�#w�"Q�%��{��<Ia���[�eonDש���E�$ɽ�*<e�bs����j��˾�[(A�Y��g��9�Y�X��ڄ�}n�iP��[P��x��F!Y�=�5G�������ל
ϙ� ��}Gδ�-����p��{��<Ia���rq��&�3�	7��ɺ2Z�'�=��>[�X��s�Q���=�����p���\	7Rn+ɽ�*<e~DN�|��]kKE��ɽ�*<eɽ�*<e��Ls\��.w"�ϕ��z	$.S����%���Hԯ��-7F:���WX46�E�Sj\�(>�g����0:��}�&gƧ)����ɽ�*<e�	S��Nd"�O��ɽ�*<e7�a'�*��wH��[�|��9f/�ɽ�*<e¼�H�4�+�T���ɽ�*<eɽ�*<eٌ���F����P�	���|v�|�ɽ�*<e��:�㗟��<�Eɽ�*<e7�a'�*����t�i��L�W��_�ܮ�	5}�ɽ�*<e��At��n4m��"�,w#ɽ�*<e�w�x�ܑ	[QI��*�Y)ꚮ��|v�|�ɽ�*<eoURqb�彵�bhF_ɽ�*<e7�a'�*��������J�p,�:��������ɽ�*<eƃ-B�ecݴ�˾�[(ɽ�*<eAn�I�ڡG��e�8���.*����v����p����x��;�	���O�8�/���%�q����d��/�z%+E�̓v�;�G��SC��Z��0�؅PSO��)��j
K�Ŏ-�ɡ���T�~��W�] �-���֬(7�{��|��5�L/%'�h���Ί�ᛢnX�0}a?K_�m�:�.��f��x�%��կ�h��Vɽ�*<ekwO�&뿃h+0��I���eJf�Ф6��4tW�,E�I������/ɽ�*<eޛfe�^C�ɽ�*<e����[�:���������G��Y��g��:���WX46�E�Sj\[S} ��I6
�,��ZQ�R�"=�Y����DФ6��4t��c@j�a��m�f�ɽ�*<e����[�:�G��cܱ��
���2ɽ�*<eɽ�*<e9����E�� ��:���c���l��yɽ�*<e}ш3�p�	[QI��(T�F(��ɽ�*<e�Xr��ɽ�*<eL�돏�㚼����|��b\	y`�ɽ�*<e�%o�������de��qw���-rvT-��P��'ɽ�*<e��}�1
��Д�٪,<Y��+�2~M3Y����A�Y��g�ݭI�ҍ��r��e�8���!���s�-ɽ�*<e��Ci��^�8��QQ>��D�\åo��Q��uɽ�*<eڵ�1G���˾�[(ɽ�*<ej&W`�)�ɽ�*<e��]{X��N��g@Z�i���!�)�49�iv (���U�n��t7�S�9P�t��^��ڄ�}n�iP��[P%��nV.�q����d��!I�2ɽ�*<eJ횈�ɽ�*<e��$]���}�M�b�eu+�'d����ɽ�*<e�1p(�G]_�,�)�q����d�3�&z	���ɽ�*<eC.Jv]0!3mk��畬�ɽ�*<e��I�v�:����p��;N{/�~:̛�#�i�e�0ɽ�*<eɽ�*<e��d�;�$��9�v��~�y���ɽ�*<eɽ�*<e-�z9�%��Nd"�O��ɽ�*<e8��T��ɽ�*<eO��B!BX��>��gʒ�D�j�)Iɽ�*<eo)���r,&�B�L^�q��9A"i�1Ų#n�lɽ�*<e�l�ᆖ���T�����	ɽ�*<eɽ�*<e���#h���U�IHomK@�Y��i;�{��5D��~��ɽ�*<e9�6���
	�P�4��0ך�������\�wɽ�*<e�ul��T�$��[�[]�wo�	h�[�j��?��8ɽ�*<e����[�:�G��c�������h���+n��ɽ�*<e9����E���=���)A�Lj}��M*71v=}ш3�p���$;���:���y��Vɽ�*<e�Xr��u:׈S�y|��5�L/%^��TfzFa+��B�\�n�I�5(�vSV��g���Ɔ��"x�N����!*�,;E��O��]�Qռ�H�!,]������Uj&��wĳ��spoz�X�}��R��Z�J���F�c�q9r�T�?:�;���A��#�P:\����u)�QX^�2���@i"M6f��������5��	"	���?��o��N�1�a�g��ۓyP������1��
O?�p٫j��"�yL�x���Ys�}�q��?Xٵ��5�,����F]�J�������	UQQ*rb�5��6��uF�p�	_�P塙@:/!M_[V�I'�
n� 70^�d�e»�-0^��,�:�	S�uP�M�zK!�g٪�'�)��F�p�	_ى�#�9�$�oWU� ����L�m�C��#��;����B�	?�gwC�N�O�lK���K)��F��P������_#Ǚ��R�����'c.�	?0-� ����Jv���,����@p~�@oH��{T��qɮ����D���,%GJ�=�rW�K�v��|�5������zWG����ʙD�0@]�����>'�6�*�q�t������ϩU�R�4�t������:Wp<!���I��d�>�r=D�9�)�Ί#|�Ӏm��!Q	s>R=��@�wG�ɽ�&���[�O�VG/"���@V��"W���à\j����f���ԝh<K��}|�?�M��\%i�������E�!��o�8���RX<���O��"P)�6�m�`�� P����Y6Z����*y����,��/�&�5K}�*���ՙ��e'�������s�SŠ��z��Qd_No���?�%6=�N����:��*D�)�=��x�Ϟep�h0����p��a!�aG���0����<`�}�)���VBm|�����N���Q�)y����:6z��Ӛ�Y���ĩ�/M����]�ͻlU��g���!5sy���tk���}Ո�,�AQ]�h�j�v���� ��B迅9DԄ�r7uo)V�&�>\���^��0*eL���J:Գ�5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�]^�h��NI���}���\ -7�G����6��_���lN�~[��>)W�j�ݗ�h��������7J�s��;H#�l�� ϑ����9�]�g�H�o*&�G܈*�\F��j�=��م�S��a���F?U��R\E���un̬���y���}�Ysn�ki`d,)�fJ������[Fv��~���OݖL�ߨ�����V��VLg-
�>^��ă�d�K^򱴃����Y�I���*qV���Բ(�~5^@�[�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�4)�}Uh����n�r�Z�}=��8����j ���T�t�g��z��Ӛ�Y���ĩ�/M����]�ͻlU����/c7K��q-TN{��UP�� �E��1�p%�F�r���4GH6�2B�T{ɽ�*<e#�\Kwz�tx�E�Bx�y��޻m�'�١�,�#S��J0�������a���F?��bb�ɽ�*<e���sz���
���Hr��a΋O��ɽ�*<ehn>��P\a��J�JqU)���������cW�ɽ�*<e>b�=�+�l��f��K�&eZ?��_^ɽ�*<eV�Q`��ɽ�*<ef��������E�\@"-��KC�F2]�J8�F2]�J8��� �z F7��2H�-��KC�F2]�J8�F2]�J8��o���ٽ�5����_k`ɽ�*<eɽ�*<e�l��m	5��Oh`�wo�	h�[ɽ�*<eɽ�*<eH�+o?�T*�D��|F2]�J8�F2]�J8�)V ٥�Dk�,���V�iYZ͆ˎ�F2]�J8�F2]�J8�T�N�:Y�?����HY3��uvfL̝g��*Kv���1Dȅ�J�_���� ��#*ɽ�*<eɽ�*<eƚ������=��c��v�5��M��̠wo�	h�[ɽ�*<e����@����xw��-����G�72L%hQQ�"^�i2���,����n����ȅ�J�_�����N���6����=�ɽ�*<e]�P�.�F� ���	/5��Oh`�wo�	h�[ɽ�*<eɽ�*<eAwo��o����] i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)XX/��m�9u	��i�\�j������rA{}u�X��V�묾/��k�P�|YZ͆ˎ���h��ܪ�f��GxN�Z廤��>,��K��<RU�"��; xX�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^��~��WFl��SC�֓�,����nQ�_�:�i	��i�\��"������ M�C�W�ڊ��4eg��*Kv�ڟ{{p��S�c�Ԋ�២x �ti�ܛ�|�F2]�J8�F2]�J8�F2]�J8�~�&T�S�p4�8��m?��I���|��N��*�D��|F2]�J8�F2]�J8�F2]�J8�F2]�J8�T�N�:Y�?�ow���FfC(h#(�:����j�=��D�z�l�v	�A)�^U�Fl��SC����a0��i�˯������L�\�ъ��7����xl'��y`���B�#�d.#W��(1�&�r��������!j�6�?�J��A)�^U�.$m�S���,����n���)-:Eߏ� ���{k����.�v�N�
�I���+W�L�i�˯����:��$ɽ�*<e
��M	�Զ���9�j�U�7v�1~@�N�A�ci�>֠�ɽ�*<e"������.��G���ʼ��9�j��sx��r��h��"��:��$ɽ�*<e��!�2X���_x�'���m��!���{v���>b�=�+�lƹ���KI�{b��D�կ��y���0	7��V��������'{�5r{#���N���h�J85'Q?�"!�����)-:E߲s}o����WVS��M`.�N�
�I���o�u�0A'�t\kz&�r��ɽ�*<eW�u���zC���2�o	����|��.E��7ۅ���|T�K�����Bj��>֠�ɽ�*<e��g ��Z.~r�/lٔ�T�2+��@�?�Vl��n��;'p�b��<���J&��Y��`�W7P�%fC�^҅��,��5K����kOe�8���)YN�
�I���+W�L�i�˯����:��$ɽ�*<eW�u���zC����xÝu�ߡ��%�h�J85'<��4ಷ��ӅT�@�N�A�ci�>֠�ɽ�*<e�s}o����WVS�.��G����G���`�wr?��pk�U4��掑~J-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�YZ͆ˎ�(�|���
4�PQ6��*�D��|F2]�J8�F2]�J8�F2]�J8�~�&T�S��.��潐��[����>"Ԇ/Q�|& ܌����sx��r��h��"��:��$ɽ�*<e8C'��h�*�U��+��Gu^ҡx�$/�%
q�s���]�[�qfy4_�I�4R������̃6!x���F�W�����[������ b��+kH�j�_�~���a�Iw�����p��@.F�rqD�h���M�>�:d�4��s$�����x��ބ~K�3������Ts�"�] ��a�ģL����h�zƈ�/w�G(j�X�S����D��m��!�'4M���/h`�7V,L��s�Ծ�/�žC���&B����7zN-���0��x�1��2��ɽ�*<e[����Eh�1�ɸ�km\9� �WY�I�F?�K���l��Yx�� �~xA�Y��g�+�r��y������F2]�J8�F2]�J8�F2]�J8�	C7��3�^��&��Z'v�}	%��)2���C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�$�䠢O)X�(�[�v���ëT�SɊ�;$�3��Q�jo	���0	7��V�IvȦ�O�9���!͌@�G��~K�3������Ts��%E��r��_� nm\9� �Wڗ�#t�sdm^S-Vd׮�8�'C�o�n�����/.��G���ʿ�Z�VwB�fC�^҅-���N�%����+��h��ܪ<��1���}��Pj��yքTX(O�_�RNa��n�	8��M/5w8�V���២x �ti�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^�M:��L���$�A����/���� ��FM�1DR���bB�깶"���u�ē;����]9]��ƅ�߼�l�G�䗅�ZC;���zP��"eI螓
JQZ�>[R #{����0��LRp����F=�y$�0�	`�EZ�wv=�z���u�@_�\($�s&6��ښ��R���C��B��1u�(���{�6ü53�v'����#�nB���I+}�p��S	��YZ͆ˎ���H����ì�Fm���W}tng
5� �����*5�_	�6���1F�����'�T �&�S�'������2�H�!����Mε�]�5�hJ�L�S��ì�Fm���W}tnA��t��4�z�t�诔Y���o���LU��t"W0�Ѵj+��njiH��gR��٘��".��U�ku5 ���"����#+8��W}tn�1U�~e&�O<ފv����%@V,.������ض��?��i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)X�A)�^U�˃�6��Rb����ĺ����Q�˃�6��Rb�i��Eta�\�H
̂�5�&K��A)�^U�Fl��SC������'Y�5a5��8���k=t\Q�w_��TE��5�l��^�ل��H�G�b��2�X C�UtVQ��5�3�4ˋ�=s*���HHs�9���h[�oɐ�c�������ٖ�H^�D����d��X	~������p���`V�f�Bɽ�*<e*��ׅ��>|
ϒ���n�78hJ����gH�6b�o�9�.\~k:��zɽ�*<e
���|H�Pk���,(nɽ�*<eɽ�*<e��ǃNICS�8�w���f6�fD�Y�WVS��!�~��y��p[����������p��ɽ�*<e5�2��5/"@+AL�Ԋ��:Y��ģL����UtVQ����O�Zl�P���;��2�r���i ;�g�D�2L.Y�����r���4GHr U�@�|-	��i�\����okRw�1w+>���֣���Fj�om��ɽ�*<e����,�4ɽ�*<eؼ��y^�ɽ�*<e�CVE�OjNx���]L�Eɽ�*<eɽ�*<e��]Z�̏�KQ��� �x8#![}|��qi��DP9���=��o��3�Yx�� �~xA�Y��gɽ�*<e�� ���{k�������v�T�d��a�:�㜋�u��F����;��2�r���iɽ�*<eɽ�*<e1��0P�7ٝGy�G��.s�x�|6f�aA�X�1�{��F2]�J8�F2]�J8�F2]�J8��� �z F7p��)Z�#N��)��0YZ͆ˎ�F2]�J8�F2]�J8�F2]�J8�F2]�J8��a��T���	ko���܌��a�W�u���zCh
r��b���9��,"�|�` � &�Wp�O]YZ͆ˎ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�)V ٥�Dk��� V
N��)��0�`�߱嚛tq�bJٕ���Ah��X�1�{��F2]�J8�F2]�J8�F2]�J8�)W���*A-�ؼ5�ob���Ow��g�.S0�Q{�5��_ʹä���:��V��9�h�J85'؛�b���-����ɽ�*<e7� �{�|�٪�Lч_%w������p��ɽ�*<e�����Q���g ��Z.��; A���]<i�HЅ�xx֔{����������?�x[���K&��`�7.\�ɽ�*<e�(�[�v���a���%SE�u)�{^��U�������p%�����h��ܪ�-�ڟ��n�78hJ��>Ѻ٤tFɽ�*<e�J4�2�|ɽ�*<eP�7ٝGy����2t����X��X��G��.s�x�����F2]�J8�F2]�J8�F2]�J8�	C7��3�^D!Qj�ǘ�0^�7�͎�$:L���![��Z�kVib�(�`O�kPNX���c+�eH���C}/�a�.�*�D��|F2]�J8�F2]�J8�F2]�J8�~�&T�S���xU�i�ӄ��k2�G�CzӇG���䜞�G4F6P�m)b��2�����=↙�vx�_1�����Ց5�^V�CVE�OjNhX���m*�f�ջ���d�r)�/U$W !��Vm0�E!ɽ�*<e��.V�+ѯ}v�>�l�4`�:�+��#yc{]�ͻlU���h�T�Rɽ�*<e�f��<j9D�m��ɽ�*<e2�s�on�e���!�f��k�2rb�-ھi��͗
ɽ�*<e$����7���ĩ��ޘ:���R)��$~)�q���������p��ɽ�*<eiT�F=U�>ɽ�*<e�ҋ\�d����#ڄɽ�*<e;�v���9�ɽ�*<eɽ�*<e� ��7��ɽ�*<e�ٱj�ꭓm�����ɽ�*<e�)�w׽�ɽ�*<eɽ�*<el2`�
��(yaf��ٿ_�6����WVS�F�W����kj�wg��ɽ�*<eɽ�*<ea��#;�Nd"�O��_�6����WVS��M`.�kj�wg��ɽ�*<eɽ�*<e�=X�Soj&��1��_�6����WVS�Awo��o��U�v�=�ɽ�*<eɽ�*<e,؏���̒�p�3>�+�{�����2�o	�o�F�-�ð�r
�z��ɽ�*<eH�7V^��uT�j�2���4�_��X�*��.�d&�������}|��qi�������/f�v"F�5�ɽ�*<e+�n�/�Gk7�����Ҵ���2�H�T��j6�C��<!�#⍈~L���V�uCMɽ�*<e���*`](0�ނT�ۄ����_g��g ��Z.3��_����KQ���ȁ`�iSwɽ�*<e~M3Y����A�Y��gu:׈S�y�:�Q�a�h.J0��	��i�\�������3X�aҥ�����L
�j0Q���'�}L�ӱ��������Uj���R�Y��ޘ:���R)��$~)�q�����b��i���sX!��Ԅ�U@�R#l�ҿ}=$�ؚ,��=cr\��}��
��<i�ܛ�|�F2]�J8�	C7��3�^��ՈW)�B&�47��i�ܛ�|�F2]�J8�	C7��3�^��~��Wɽ�*<eɽ�*<e>"��;a��yl2���ɽ�*<eɽ�*<e`ύ���#�k�:��X�1�{��F2]�J8�����q��2������J�e�m��8[�5����fF2]�J8�$�䠢O)X�5��M���>���6��ɽ�*<e~4�R�T���5�W���.�^<�
:�ɽ�*<e�&�|�D� ���	/5��Oh`�wo�	h�[ɽ�*<e��!�2X����]��5�5��M���>���6��ɽ�*<e��)����;�&���i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�)V ٥�Dk�JC��������>-VV :�>�51�yƾ*�D��|F2]�J8�F2]�J8�F2]�J8�>s�^�Ym�1 ���j���@n��(�6�g��IϜ&q�t�	��Ę�:4;�hO�<���J&̊��5�0;���ic��ݤ��:4;�hO�<���J& 칽�y������[!����q��`6o��f��<ߔ��:��$�L��g}���%�����>��
��`6o��f��<ߔ��:��$�L��g}���%�����4h�6�`6o��f��<ߔ��:��$���&U=�<M�h
��Y����^	>E�I����������4h�6�`6o��f��<ߔ��&�ӱ��k�/�wM�h
��Y����^	>E�I��������Z�7��4h�6�yr���wٕI�+2I��!&)�@���0�.������;�*(�h�A+D��R�×_� �)y��C4��;�Q���<��%��ݝ{w91��?���,�`��� r��B�@��DLno{Q��+���\	jG{{�h��xt�%��}<��B�#~���c5.Q_J�=�ȭ6V�;4����z8����S��z+t6��y��4��<*�o�A[��,��)=�-h?>4�DLno{Q��+���\�S���FC��]�����������4Cxl$5Q�I��*>J
�ڝ�1�V�\,��j����s�)���_:�HS����ۖ�hh�*��.�d&�	jG{{�h����?5/���05N) ��񁯶g}���Ps*�^�j̇�E��5�l�0�ނT��\�ǋS��<�Q�E3#:%� 2]�������F2]�J8�F2]�J8�F2]�J8�$�䠢O)X�����)0��>v���E�J�����u��S�e�m��8[�5����fF2]�J8�F2]�J8�F2]�J8�T�N�:Y�?��טZ��9˖�����X#�����;��y� r�Km���¨��q��v{�븽�Z�Q�_�q����O�(��hܦU�*�J喌(��0�X~_�L��I`�a 4�T� �' �.���C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�*"T��v�
���ji���f�<�~��ݝ{wAwo��o�x�[���p�v^����|��.�}����u�9ݓN��s�KYyع]�0��H�m?�GE�'^����]���W/�f1�̕������,b��x E�3�>�����u^ҡx�$�~'d�5}�R�ʹXr�	e���)Cm��Fo�l���2+��V,L��s�Ԧ�yB9�O���U�8�s���2+��ɽ�*<eV,L��s����C���������>P:j���"��-G��g�f�P+txP:j���"@�3aăP��8t����Yr5�ŕI�(^�GJ��a��ɽ�*<ex��*��~��h������?R�0�"��*���<��lk�/�w��V��RvS+ё@{���W?t�<�Q�E4�+����ɽ�*<e�@A����+�r��y������F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S���s콻��ۭ�����n��ZJ�d�����:�3���"��; xt��f+�v\����
D��˶\Ȩy.1"^�)?��w@��*���p�?��x#���G����tt'G���XBg!����M��Y���j���S�tYA{}u�X�y.1"^�<T���9��ė0��R��:���h�QU��c\���e*�����W�݋5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�u^ҡx�$f:@��L��CVE�OjNx���]L�Eɽ�*<e}��黯p�,�3�0+CǺ�Q���\�e�=l�^a�M�#�C��q����ow��{8[v��c��޸���s����ɽ�*<e
���|H�P�vԻ��;�\�e�=l�/(� U�A��K��k��W-��͡�}Gδ�-]��ʣ�G�H/l��_)�:S�c�T�A�Em�\f���}\��hߡ�8|�t*lC60H��r�dZɽ�*<e��8t���՟�>U�G����R_�f	.�W��t�]��#�ɽ�*<ex��*��~�������ɽ�*<e�ngF��U e1#��A��K������p��ɽ�*<eO�
����~�|�)ݑ0�՜�ıU쏘����K�^ׯ0�ɽ�*<eɽ�*<e�\�e�=l�/(� U�T��T����f��Ƨ�0��+#�{T��%z�@�(�=ā~�XT'�P�.U�[�x�l�MȁUN�\�mI�V�A�/�l<~OX����B�8�H`���@r���28��&�������p��O�
�����GbY�%�����p��ɽ�*<e�`V�f�Bɽ�*<eɽ�*<e�������f&�Rk��ɽ�*<eɽ�*<e$-t�O��E��o��ɽ�*<e'$��R��e�����kV�'$��R��e%�̋]��ɽ�*<eV,L��s��A얺��Bɽ�*<eɽ�*<e�#`LL�%�oX�t�����h�ɽ�*<eɽ�*<e�)����>#	f�
�+���cP�Tɽ�*<e��8t������p��2D��B�i�ܛ�|�F2]�J8�$�䠢O)Xv8�����0�`�+g�Qt�C��ଡ଼�F2]�J8�F2]�J8����4T!����tQ<[��"��	t�nQ�ɽ�*<ewRۣB���d��-QJɽ�*<e���npX�����p��]�P�.�F����P�ɽ�*<eE	U�`�x����&�����@���ݝ{wAwo��o�o���l�L�T�2+��@$�sA���[��v��/[3۷_=E��Rx�����y���yO]�&��I���R��A|`�$������kȡ�B,ŭ_
j�����ͬT$OeMS���s�C�罤�9.�f�i����
D��H7����{�ƥUuh��V�g5D�l��9q�X�:׮�5:��KL����z�>�4[���{u�^ק��}�{�ʘ��SD!��Ю���0�V�٦�����2���X�����wD`֡��y����"�m���F^��`���#H����^'�2����:W�0s�����S�_>gN�-�:'��$+���G(����^Le�0�[��z����jcbb_�B�,��y8f���B6Km���'�5uEq_�<|7.���|N;X�^�I�[\o|�o�����|"ÝW}�utiO����+�%�Q)=d���E,��h��DZ�x���F\��w�0��8w���c�Y�l�%�tB�*��� �&&s�:v3�9?k����Q������L�����p�N_�qe�
��>̊��%�
�T���k���g���*�F/��q+�\��$|?G��a�G�x�D�9ϑm�eQ���9*Q����� P�7+��$-���G[�z�A��ie�\#�_Hc����'d����uC)�E���Q�0)Dm*
kma��ݑ�`��N��X5/�)I�|��o9�H[��UF�n]h�^�o��p����=����+P
���(�5;B�W��M��v��E�`�w$�P��j�:�mheˣ��:��?Dg,2ms����{Ue#T&�ީ�q�� B����ڴ���;������kȡ�B,ŭ_
j�����ͬT$OeMS���s�C�罤�9聯�v!�������k{��Ty}�zj�"��0��U��j )���.s���2D��%_�y��N�[\��NT��>n.r�P�S��И]h����,��D�se��L���Ӡ��B:l��9q؟��?��6\F�߉�}3z�s"�!6���f����!Lؒ&�bL�.��. ����lB��,zyj���0_��A�\��B�N��%졖*��j)?��(a�����@��$�G#�ӵI�0��#Ҟ�s�-I@>������BP�\_�0'���I"ʈ�W�rB�������i0aXK��2��H����D���i�6 ��Z�)a��\ `L����B)JǴ��	ĭ��n�W���\?�R�?3�h0)�E�Z��(w
�7`�	�6�����C��F���Y��U��>��M���2�أ���Q������L�����p�N_�qe�
��>̊��%�
�T���k���g���*�F/��q+�\��$|?G��a�G�x�D�9ϑm�eQ���9*Q����� P�7+��$-���G[�z�A��ie�\#�_Hc����'d����uC)�E���Q�0)Dm*
kma���t�jp�]$u�	8'��v�eMV�z�U܉����4�=z��F		DAu��6YhzoC-x�i���
V�r&A�V�6�.j���|R��Ǥ_�|�P��L���Xj��)�*��e/6�5��0�K(8 �%D\������A���UJ�l�t�p,|4�^,e�I��ހVh��S�zC��YB�gN2E[5���ԉ[��Q�)y����:6ݑ��/�׸s7��s�����Ɯ�h�Z��g)/x�*B��0�ѡlv���tk���I���v�D�t*�gc�꺉�@jB��Z�!�W�/�CQ,^�п�cψ5����4���m.����c���5\�YuG���0��Jf�x�\("��	�wR"]�ͻlU���(�����iP�8��J�=�B9�+�й���M,�Q�.#��K?��MT�6��_S�%���t��*����S7Wcq*�R#l�TB��G�o"	9��Fgɽ�*<e �����2}FAt+=�.��ԟ��6�����H�T��qɽ�*<e{*o��^]��������J�^̍�g�z}v�?�vɽ�*<e��b7A�:2}FAt+=�.��ԟ��:9y����B�p�?�ɽ�*<e����J����DF��t!;��[?�����Njɽ�*<er���4GH�"��bdA�p~rև��h����hǳ�o�ɽ�*<e�����g�Hq-TN{��U�R�.���eif���ɽ�*<eɽ�*<e�2a	;!7#]���������ݰw�x��\t{Đ��-��!�G��b7A�:�N�]g1,�Q�k��/�
��
���t�U�Y "�t��{d�.{d��jI-ɩM,�Q�.#��K?��MT`q��Z�@T�R��n��*��s�� 7���]���������ݰw�xo���R�-�	F��ݏ���f�W��1���Q�k��/�
��
�����$S�ƾɽ�*<et�I=1��M,�Q�.#��K?��MTHk�K{�ԵL	��D2��*��z�;!UF�R#l�h"����z���6sy�ɽ�*<e�q�҇�{�2}FAt+=�.��ԟ��� Nb '�B��K�ɽ�*<e��cb|���DF��t!;��[?��$(�dH�T��qr���4GH�!�\b�ڬ�p~rև6%�p=��4�d���ɽ�*<e<*^�i�q-TN{��U�R�.���� ����~��0�K��ɽ�*<e�N��&���]������ˣO_���!L�E�I6�L	��D2��b7A�:�/?@؄�-�Q�k��/�-�]�x�{ ���(5%ɽ�*<e�et�}-M,�Q�.#��K?��MTJ�k2����J��V2f��*��.���̘Hq�R#l���wwU���C �7� �G?�L���m�x!��2}FAt+=�.��ԟ��tV��^���>�A*��O2�9�L>0�>��FT��DF��t!;��[?�sN��8H��!���pXRY�Ȝ4�Jf�+���p~rև6%�p=�O�;8W�fL	��D2h	Ӎu2�q-TN{��U�R�.�;��:^��Z���Kzaɽ�*<eX�n"�.��]�������?|�'�v�<l]j^a5k:e�."z;� v��S
���j�o��Q�k��/���0��Y"�����Q��V��~��X��K%��M,�Q�.#�1�e�xHB�P�.a7)�ɽ�*<e��*��2��ȭ�R#l�5jF�߅��!?�)�ɽ�*<eQi�{Ѩa ` ��Lg�+�4 ��p~rև����/�WiUo�	8��~e��H�`_ɽ�*<e��#�Nz��=���øxQ@Q�;]2���U��DF��t�N\�C¦P�.a7)��/r	� �6������D���ts��T���6�e��M��p~rև�)��@=����L�N��K�N.��O��DF��t!;��[?�dC�r��w; ^ӭ+P��FB^���)$�zsK''oB� ` ��Lg���p��������[��J�й���M,�Q�.#�k��ot4�hɔ��|BjT;�9��n�����M,�Q�.#�q�����^�V�ɝ�����-�~�F� Xv1�0;M,�Q�.#��W*͓MfKˍʔ��	kU�f�Z"-w��-M,�Q�.#��W*͓M\�j׸'��^H"-w��-�un����_�Fe@�[ݧ/��й���M,�Q�.#��d��\V�v׿��b�-�]�x�f�5~��r:9y����?K��qq-TN{��U��rb�����b2ޏ��O��%Ȁ�un����44�f�K�x�zW�ɢ�.�֏O��hb;��?$x�U �qO$�a�Ow�6N�]��&�]�� �pz`�<49&n���o�t��p~rևu�����j�;��T��ɊF;z5����_k`ɽ�*<eɽ�*<e���r�<H�ڸ��P��B�a�h�ɽ�*<eɽ�*<e`ύ���# ` ��Lg�Q��t�/�F�W�)7��NVUl��؈gVy �v-�h�!��qj)�0�V-�����B�Ja�f�ٱ��
���2��
�a��;� �:��;�X�>��]WOao@	�;0�头�˾�[(��
�a��;� �:'�`}0����)-:E߁+��>@���b\	y`���
�a��.�^<�
:�ɽ�*<eɽ�*<e�������J\]�n�z��e�j}}��ǀ�Z�|�CEP�W`c-�b��"/���?��H�ڸ��P��B�a�h�ɽ�*<eɽ�*<e
Q���Ȃ��9����	��y�i�q�k�אɽ�*<eɽ�*<e8;��4RȌ)squ�`�)����N����1{bhA*}|��r8�1���E�Ȯ�^q.J1ȅ�J�_�\�I;���ɽ�*<eɽ�*<e�Ja�f�ٿ�P�6;7}q�cW����5��M��̠wo�	h�[ɽ�*<eɽ�*<e����Bt@��K�,���Zr%�����B�a�h�ɽ�*<eɽ�*<eEC�[L���%+�mYr`����&��S�Ƃ��ɽ�*<e��*?�5_+�v�i}�"�a->�d�wo�	h�[ɽ�*<eɽ�*<exP,v�L{���V��'x�|���C}�/��c�y� U����e��a���D9$u�R}c��̠!7Ni�9�@q�w28բ7��7���G�U�E;��]��3�w�;�o0w�7����&P0��GA��L��ְR�	_��%��3\�!ќ����,����P�C����е���09ӵ5��L�f�����ȶ�:j��,���?��-No�bg��@<�i"��q��WY��¾ߝ)���{�_bD`9�8&�%�ޅ�8��\#����r��{�t����s��v���[Dް�F���W<:K��cl�V��C��s�ߢmq�\F���P�V?�������7�5��M��̠wo�	h�[ɽ�*<eɽ�*<e�B֊ ��f+��c���
�a��.�^<�
:�ɽ�*<eɽ�*<e�5��[1g�R�a�G��̸B������f�U���6?���:�ɽ�*<eɽ�*<eG�k`>-:��PO�K����<���^:{��ſ5����_k`ɽ�*<eɽ�*<eG�k`>-:ÙEǛ'�s^q&/h.hX�����2�R9��ǔ�[$As��d��q���EU:�h�H�yl2�����(SM+T$J�{7D���)-:E߭�*�M���H�KV��iI��~��Wɽ�*<eɽ�*<eɽ�*<e�5�MP��=��c��v��~��Wɽ�*<eɽ�*<eɽ�*<e�5�MP�⠽���d<�s��7Z��~��Wɽ�*<eɽ�*<eɽ�*<e�5�MP��˃�6��Rb=LU[$"�eF9YH,ɽ�*<eɽ�*<e����2��.����Ar{@ �P�G
�CL�;Qi��e��E�JQ�.x��82��5�/���J�����Xĥ�\#����r��i���K�9�xQ�����3��Z4qP�:g0��4sN��8H��&�ZC�$R�5��M���*����/��ڗ��`���)-:E�����M�L�����`�yN�F�8I����N���ɽ�*<eɽ�*<evS+ё@�[V�`��zǙ�7����k�L�\�I;���ɽ�*<eɽ�*<e�f�P+tx�X�Bh�W.����T�3dHL�`I\�ʇ5dL3\�!ќ������S����m�C�<��cD}��G�P�!oI���ܔK�"J����vS+ё@�[V�`���>��h�
ȅ�J�_�\�I;���ɽ�*<eɽ�*<e�f�P+tx�X�Bh�W�	�y{I�7���k�L��eF9YH,ɽ�*<eɽ�*<e�f�P+tx�X�Bh�W��.����AMҼ��>i\�I;���ɽ�*<eɽ�*<e�f�P+tx�X�Bh�WJ8�-�3!Lr�5"�O��
�CL�;Q5�yj�N�d&f��E�*vU�L��GEU:�h�H�5��M��̠wo�	h�[ɽ�*<eɽ�*<ey�1�+·��t��.�^<�
:�ɽ�*<eɽ�*<eĳ���|w�ac]8���}��G�P�!�h���*b�mq�\F:j���+�@��4�(y�yl2�����h�����V��H�f�������B"�ހ�l�,H_\�I;���ɽ�*<eɽ�*<eiԙ�&�Vb"�#F��87U*���g�yl2���ɽ�*<eɽ�*<eɽ�*<e��P��l����F���C}�/��c�C*	�����Iܑ�LZ����`�g�v���e[Dް�F��~��Wɽ�*<eɽ�*<eɽ�*<e(��ʸGଟ�
�a���f�[>���ɽ�*<eɽ�*<eB�+��������k�L��Kn�:O���B�$J�{7D�+M֏��_H�KV��iI���W<:Kɽ�*<eɽ�*<eɽ�*<ew荦xy�cV8��+ Z��
�a��.�^<�
:�ɽ�*<eɽ�*<ef&��7��f�K�am@��k�h�������F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)X�����j�Ԩ[��d�V��{|r[�i��E�%�r�-?��@y���V�5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^����2�f3�I�^S*���������ظ��~��W�v��Jݍ���!D��'ί�|ޞ<�	�`�lpŌ3�6K��V,L��s�Ծ�/�žCq)�_��C
�V[�?��=��5Fa�Jg1�4�b�z�atG����ie� t�e ��:��%�������.t���90��Z[����x��F�Y>u���kɽ�*<e9Ӧ�^�q}��̫'ɽ�*<e1��0����,�4=�������)��՞z��߿X�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8������MP�J����y uA�6[���l�VUQ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S�=c@�LT�G�di!�4�^*�����ԡ�ZPZ�-��K#��]?@���Hs���JYw�8�r�rz��bm��L2��/r	� �:9y����HQ���y{`is3Z˨��ҮE=c@�LT�O�W��̴S˝�#F4��ԡ�ZPHk�K{�Ե�D���tsY;������	q�ho?nr����˩�En��G���]iLC���M7z����9���=}�J�vMWK5�ޭ 	q�ho?nr�����Va�I`!�◜��y�>4�*��@L�E�I6��D���tsΔ��B������ҮE=c@�LT4���v{}��ჭ�u�l��U�Oa͓܌����B��!cQcr�j�����2�O��BB	Zݪ+i��c}�&
Z���dZ�D6%�p=�O�;8W�f�D���ts�����Q��Y��o����JYw�8�r�rz���(����vr�0��@�9�P���95�c�V:��=�
�nr�����`��ʵ���ȃ�?i\C����D�/�	��l����L�N����5�=c@�LT4���v{}�f"��w�>���.��J�)�����A�ֻ�mԳ�l�VUQ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S����=��g�Qt������F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q��1q5	R-u��<,�A?2v��<uM�Dl�7�����с���-p��V�����B���L��J���1Ѡ�{v���j)�0�V-�����Bt Եp��rw���F�v�hR/�͢mq�\F�%,!u�r�	:��v3h"J��D(�R��-�S�Ƃ���D�r�"�����сɽ�*<eɽ�*<e����Ǣ���O�F��:����Zɽ�*<e:j���+�P���B�'�=�3��&ꬶ�Rɽ�*<e�0{�I����՝��0s9�>��b�zN�����ɽ�*<e �jv�5�=da���_�'�=�3����,g=%�1�8���g��;i�m˧�s��'�=�3���%�p-�djJu����<�e�/�{T_��ë��������V��P�����|�kG�qТ�j��ԩ����;q����n�zN�����ɽ�*<e �jv�5�=���W��K-��'D���A)�^U�ɽ�*<eɽ�*<e��3�y��X������A)�^U�ɽ�*<eɽ�*<e���8o��%#�&�u��I@T��Z������ɽ�*<e��|s9�,L��b�!ȓ%�����zN�����ɽ�*<e���Af/�(��i͛���0�RKD�vQFɽ�*<eɽ�*<eª઱ތ��I��ʟxҦ �l�C�'�=�3��&ꬶ�Rɽ�*<eT`�(O��2#_w����;
E7���������M�d2�i�(�A��q��Uk�g�uQ�{U�y".�!�M��*���e|X���XgM�] ��?Hs�	�j(�d�A�S�Te�Mf	h��]L�/>aŞ���0��� �H,��~
�H�8�c>����:9y�����2v��AS�����Q��R&�'�Dɽ�*<e���N�SVMr2����0:{�y�i�USm��]�Go>Q�צo}��Pj��8��ם�5`��)���aW�b9t�ؠ0v3>"CA��e���l�O�psc�w5��*�(�[�v�����h����I��c�eŞw�=px����`q��Z�7U�'R��(�[�v��25�ΆQWk�HZ�c�eŞw�=px�������������M����}��Pj �e�g0Nd"�O���aW�b9t�ؠ0v3>u���|��G�@<O�G3h��]L���-c�kɽ�*<eH,��~{��\�jb��{�?��e�>��9�����Ym}��Pj|v�cɽ�*<e�aW�b9t�ؠ0v3>�$(�dOYD��ˣ��Ez`r��q�Qy[�^N��k��ő���s��l�u�I%�F������L�"�YZ���x;< ���:94��x��
}��Pj��:�JXL�T�F*=��aW�b9t�ؠ0v3>�P��Tiu8}�̴�P��Ti)�8	�q�g�����Q�I2��)��|T_ӷ����N�SF� tђ�.�w <>k�qH4^�v������Q���TU��}��Pj�O�@cn㗟��<�E�aW�b9t�ؠ0v3>��~�1�7
�X��dR�J]{�ΓJL;kAt���
+7}��!�O���=?э�@�R����,�"_VZ{G�{�
��\���(0.�溃Z)m���e�u_��F��F�e���Qq���,)%R�i?21Q�W��P�{�[�#t{u�$p8�2E-�)��#U�$^۱�j}0-�2���:WY��n�Av�'�B��w�Z<�{n�&�i�֧�d���;%�s�Jq��Y]SҀ����e!Ju-�!�J�`���m�)[�% ~����j�(���ft�G4Ġ����`�K�"��ck#*H.�F%��\�Ϻ�x����F�K"����Y����ƭ��wf*�.�P��A)�^U��������n�����m)v��V"��`~!h���7�E�"�w��tn�[9���cs�px�����IuW��Od#��1���F�2'H?��R��$�,4"5˭�����������L\�`�P�J��w��.�����с:�)�A�08�bB�[�Ͽ()zӺ_g�=Dٛqוۏ�.�E>2�<U���	��wF��2�,��6�/�9FO��G;ϼ^�� ꫂEޘ�-���Ծ��#��V�C�2w��Z[߷�J��'�=�3���|�T�C�p7���_�8����		%2�>��1���L��P�0��W�d���y�j�(�h2��M2|B�7ׅ�|�7}��K�am@����:M����P?���ݚwH��(yv����$ӟ�V��\K$%�,�	/ؠ���'���
�ӴW���Z�d�e�:^(X;��:`�[�8�'���p0����сZ4�Q*#9?��{�h?e��NIl�N��Q��
ugkbֿ�S4�ڹ��lΔ��B���bl�acui+�ꤡQ�`w��g�.S��}Gδ�-�QF��V��:��k���DC0-�'zxrF�h�(�Vպ�ͫ@LȪӖ2}�nQ=͗�O���-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�M��X�{���h�<���\$�� ���3E��HdAI,�FP�X��D��)&�"<�tL�Ba�O�)�\�zq �����p����`,��T�VJUT���j;tZ��k����%��+<�+`��r�8�m������/�űё�L���o�-M+ɽ�*<ezb�"O�a�Vz`�N�:��G�1�&��Jr�Wy�~�(��V�?U���3�B 8raɽ�*<ez��B �
E
�P2t�s�U�F4_ǔ�m��R�U��6~JV5	� f��V3�����p���㕋<rt�t|o[��H���/�k��|"ÝW5�/�S�ҏi�$:3���\$�� �N�f�	�e����n��r�o+\��&�VJUT���)!)gP\�@�y��F�g]�VPϛ<,�dBh]��< f��V3��}���u	|�5%��Ż.=գ`,C<.�ދ����������n��rW�񌷸:��3�-��i�U�fw���H�~�����%D�]_�����OQ1�� ��1A:���ɽ�*<e�&�=A����Gn=�(�v�e�ԝ��E�QRH�l1â,6|����=A:>�m�V�]�'"�79ɽ�*<e�����|W�meju��*F���r}�y�:�#�Z\#�-C�����y>��XG�GMm
\��L�ɽ�*<eT�M����24��!�굲(�x��m	:�R��.L��,QR^!*��|ģ`[B����d�v�����AI(�w������p���G����G�QJ	�i�4�c�C�����rɇo�G*�T�tȈX�?nC�����/�űё�L ����[Y���o�f���^�?���2DC?�Y3�~�`�/�HY �����Ǫ�^��vD��9�����b��.I�9�PW�#���;v�a�GO��}�w��_Qgs/�űё�Ll�|���N�|ۈ�;�Gla�Jp����/m/b��}F�\ɽ�*<e�%i��I�I��u@(�o[��/��$��E���`�
��q��G������Vɽ�*<e�����F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S�����p��}��PjƓ�pp�\�鬧�N�׈���g�ÙEǛ'��\DԷ��JkwO�&뿃��^���۵��g���>M@���a���9�����z6%���TJ�3��&ن�o_�Iet���
+7���1b7�&Nꊓ�HL�"۠����GB���,�6}:&9%a��ە����7��h��Rj���ɽ�*<eihC�^8[��(��t���cU���)*�Qy*P,hc�Mdu�h��q�i�K���^ưVx}��_������n��g9�� <�t-*�����p��}��PjƓ�pp�\�鬧�N��6f��C
�V[��h�<���\$�� m��-C�C�.�(�.����;�V�`��ɽ�*<eh��]L�;���7d/��c#U��9�����z6%���TJ�3��&�4�b�z�a�+�r��y�Q���'�}�ٔ^qt����g�H�D�V!f4V�ɝ�����-�~�F?�9���K�9�9�d��PtD��v�s�ɀ�>�8��d�f��D)�Y6J|X���%\	V�6�}��Pj�*�^���lQ���=�1�pt�6����d�՗�*3ZC�q�:�Uez�|��`�$��������\�ռ]��h(|�%#�&�u���`�7.\�����Q��5f��˵&�ӂ[u�{����/�;� �D�w�,�o,�����(�[�v����6u���}�sL9?�Ep�b]�gD^t=�&E�i�}�x��r�֏��9��&�[B�8/�2!�ӣ��$n@��L,�|��b��!��\���Hb;g�v�s�ɀ�>�8��d��btX�８��%j(��Î�HX^|�ݲW��;n������o�)'A��;�����)��h�(�[�v����6u���g@]l�I	�p�b]�gD^t=�&E�i�}�x���j�8]��O�j�<��{�
�'�r��72^o��t���y�P�(�[�v����6u���}�sL9?�Ep�b]�gD^t=�&EژM*昜n �e�g0���T䝎L��Ԝ��5!��s5�;Ga �>Lp�G&DQ�^B%�(��Î�HX�Iҗ��nL��b�!r�9d�x.���\!�����^/a�7{|��8}T�P�ԧ��Fn�p�-W_xZ��C�}��Pj�v�s�ɀkç�$|i7ǉ7ҡ=M�%���K�:�[��P�X��X���l�VUQ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�HE��޻'���'�T�Z��:�^4�M�(�bJRܿ�Y��4�*29���Ι4{yP���5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)X�c�|ItȰ�4����y
���� i��1ي�b������J�76Z��p��P�:2]�6鯷����`"�Q��B˟�����p��%��jHi�S�"����*�#����o"s86��{%:�?l���5!o_��^^�V��6Gum�?*�����&)��n��T݇í�ĭ�U��c$���
����뙙_	=(���U>�,�x�u�o��1و�d�Q���TB�'�~��5�w>�8F�]>�F��:�o��\��?�n��߉�.�CN],�'�]�m1��@o�c^��� k�n�� +0iT�̰^�*+�mk����͹ �_d9�p1H|�'ࠁVk�'r-�c�*�/��0U�|mD=R���Y�_;�\ `L���N���t�E��'�MS>'�Vї�$te���n��좋��N���� u`�i��Xc��iA'-{�>�{u NEzʠu8Vr�ǖ .�����#�"Ӆ�g�v�-�t�؂&t��b6Ԝ�,2�����gł��*N���D|.��T��R۳R�>j���A�u���4t%,��{�	?�^2�՚8��%g!FBRi���D-52II�.䫓�-��b ��I[VfW�a�`����M��_D7��h�¾�Z=-�ݞ�Խ��X�BE�����f����UH�Xzd��7?�Z�'����!�O�
����V����H�oM�1�y<1l�XiI�{��2j#��Δm�������p��}��Pj�V��S�*�іyo����R&�'�D�^��+���<�8�֌i�B�k-�^��g�7����m�u�?~֒��a�ߔG�=����<��ݭd��PtD��m��d���
���2�ߔG�=���(�[�v���s���0��z����Q�H�6$���ߔG�=��3��֪��	D�ܣ{U��m����?�s��Д�٪,Ӑ��4�&4�OI�:q�Qy[�^N�����^|��]`��(c+~����{�>p�|���FS��J�^k�?���_N��^�Ȫ��d�����N�"J��6?��f��?v!��)�5`��)���+z%~�O���D��"���8���`9r��aN�#
@`��w�N���]�	�Ϡ��)1�،Hߜ��'��ø�ڠvs֓'��4JJ�Л�t.X&�@��N�O���K_�[�'-qR�o��}tj�� ry�2��I��F��,g��/��b�?�GaӔ��ҐX��w��Z� �Zk�b�xk��<4$1�:◥�o��9sW�ɭ���U�E�����W_�G"��5{ �3=HǎXJ�76Z��p��Ѻ�/��ZK�;�V���4����,��,�;�Z>/~���C�)��w^�e�kny�2�PO�l�c��I��V1��ܽ�Sp$P��Uۭ��H��3��*����U&'{]L�D����y�%Q��f>�N �A�gǋڇ�'T?^=�VC�oʄ��Ck�,�G��Xùo,Mh���/���k����I��ܨL4b�ްL+�\ݣ�ӔO���MG>���d]�@��pz0�Y�Ạ�~L���U��;"�1F�X�Pyv��*���w��>��Z��ĺ���~��O�^ZY����՝����돷��Y�u�}��ޱѨ��t[�����Q���s<%��`-<2N5}��XUq��ܶ7��R1�c�9U�H<̅9��4S�\��{��̠o�����I���j
(W8%�0܃DmaXƻ�2��|
�V�|x�w~0>T���;�X����E��L"�~��Ӏ��mф����\m�l����X��FQ��(�A�c������d�}_�3��$S��Ak委f�*�i�� �7�7�Om��������{��\K$%���	��o�t�%�j���^�hq>Qm�D�U��eNܚ�d�Ŷ��T/�x���LI(�[�eonD��0��t!h�a�$�ou�d���t�Q S-E�c~:s�m]��ȋ~`�}:TM�E�I6���,����n�m����P�/�k���	A��ŏ=����V��+�j�+��������eR>��h�ɽ�*<e}��Pj��E�1��kv�S���)�|C�xE<�=mArА�\��{��̠o���a_��k������p����+&:���^04%�F�}3���~��ڒ�ɽ�*<e;�\u�U������4ƕo�Z���uȔ
��pu:׈S�y|��5�L/%}�tؤ�l����������D�\åH=>���JU�I+��j�8]����P�*�J�EL�cm��H��1sw}��@뾢� 4kZ���6�/�9FO��G;Ϣ�>U����\�e�=lS?�1e@�۱�����tQ�onv>�v���I�q�)� �)X �jv�5�=��4�B���%�!z�Q�onv>�v���I�q�A�Y��g�+�r��y�Q���'�}�ٔ^qt��@�i�zr(HU�Q`-<2N5}��XUq�Ά��#��@?��R���	U6GI!��@A����6��U���@�i�z��{�\w6�`-<2N5}��XUq�Ά��#��@�OCs�Ћ�e�F�g��5�h��q��֎*b~�*����n4C�!ʑ���,�IM�+�I���0��>�������h�fd�	m�LC��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�:-ɭ�*<CF��͸��V��[! iZ����`��!9*6rP���Uq� ���}(H"h�b&�� }�I�Z|�!�SY��<�0���ip^6�HdAI,�FP�_�`��'����Tү���HԈ���$�1�du7L:լ��~�*(�6����օ����� T�u�R}c��:#�̐*��=��<���/sXI��XR%�-��h�'yO�x�+%�߾�>&�dO	�0DN��1F7�C��\�c+��I���>�~彄W���^�IoEν�ڇ
�܎[2A���U�ָi�Z$)�]��d�|�L��5:U<���=L�s�biL�.`�d �|w��@?}�Č&���V!�F���t����jܞ��VCø��A���9ަbq<Z�Gԍ"ώ**����7�#�g;I���)TK�o�NQ�sK�R,�FZ�������t����8 j-�ޡϴ��ܳCǢ�klc�+�3�g���fr2���G[�t��NxL �?ղ
�L	��F�������R���M�NxL �?.v*M�K�\��ڬ�t0w�C=[���V��Tf���9TI��~-y7�6DL����z�IYLy�0�X���p)2���@�h2uv<�WV
v��
���jiЁ[V�`���S�)n%�U9����2X0u0�pM�>�~1����buE �}�S�axVX�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�&���y���s��������ڔy)i��y1�d�d�Ɛ����r�~}M��W� $�Zp3�E��.Ȗ��@� ��0�)�֣�?����m�6��9��ڇ
�܎[,���7I\�:L7�B�e�+��U�1?�	>E�S� o׿���i�NF�X���kEry���k���!]�4u�?赑X�r@�2<b�]łB�w����#<�}�AͰ74dv�ڇ
�܎[�V�²z<ru�R}c��kOwԫ��蚊�?ȴ倠�.�Z�N�����D�h�r�<�����5`��)���R���n�m^.��S-��^�,m^$cI80���h&� ͞����E�Ի��(�Ǭ.ɑ�0��~�~&w@���m4��(�%����#�_v�jm�}y��������B��{�4���~FKV�L�ߨ���`
΁����"���A�R0;��L�S��ō0�/�����m���SN�kI�?:s�v�i}�"�EϬ�^[��z�u�!�F�d-��寢�2Sn섮@��PE��+*#��ّC�ho��9���l��K�֋3̆�B�_.�M��W� $��j���t��f.��d����lZ�����9���瓓!X�ω|� z(��/3��V�/�C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S��A)�^U�(Sg1��կ1n�W�o��H�*I�}��Pj�����Voցt+�5%�V�²z<r9|��P)U�w:����S�E �����6�/�9FO��G;��鯶Ŧ%��J�w>����B���ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�/���%�&�R������=��Z	��Ͳ��^5�� �	(Sg1����K�am@���P�,(`�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e=;+��.��d=MK(�b�sN��8H�����zxᪧN�JFi�2�5�}�Ň��O#�!��@A���H�Hk��Ne�����%��k���a���D9$ý	f��)t7�8Ҍ���#�_v�H������R0;��L+�ʲ�R��Z�s�H����_�7���X� 9�^�Y�@���y�ɾXe�gc�8�g7�-�?�d��V�P���T���s�D{�.V���6��z�<F�	j�֏�d��+
�i���<���^eZ��K�����֟n�j�T�FU)���7a��}�Nj�$9t��xl�	u�R}c���9ަbq<���>��~��V�²z<r�Ұ���ɾXe�g�u�z�|em�n��U�H�f��F��V;*'76Ǳ� W�@Q�;����v���O�t4�.�2~ ]:Z�NW��Mdu�h��/! �f5��#�9<IcX�ל<�����B� __�DȁA�>�6ͤ�PFw�ݼw��kjJi&'��t/:�P���-0Kl�c�"�=�z���b2�R9���V}ڗd9�^5:%�|@�������^5�����9�7a*/����z��<�?�9����{Q�! ~�$��A)�^U����YuI��P=�{"|`�_w�A)�^U�s�ڢ>��OFަki4 .pK�/�M��n�
q95�c�V6�΂��4
�D��ت0���o�P���P�m�m�ϙgS��^�hq>Q�&w�z2���Z&2��[��K��\���c\(�(�[�v��w~b��虁U��A�w��*�p�. ��ޭ�\�7m擟��"`�˨ƿ��;�X�>��]WOao���T�
�1����w�V�!GA>��E�����}$�$`����Z���u��k���>;ǄN���E,���T��)\���J�w����#`x%��o`.�E���cC�?��R���
�\۾��eO�(�Gj��q��y�[��)Z��
���ji� ��w���&��N���|C�xE<���&�;��8�T�ȷ#5�|vk����#�>���`܋f�~��˃�6��Rb�&;���g�M�9�mćX�V�?`����M4#�$���$t�_rw���+��]��#�p�xN�Ux��I.d
�ԓ�M2|B�7��>��R�ɽ�*<eɽ�*<eɽ�*<e��ײz�'��XUq��;�4ǁ�ǉ�T�2+��@�(�[�v��L��KN�Z�j"�nm�B���uVC�<"G5�td'-�f��ݬ�����Q����P�V?8����		%�����ofQ6���V8��+ ZYBDt�@$��[��Ƹx���]L�E7�����\���}G�5�28�W�� �ʻֻ�CL�!&�����y���|"ÝW\#����r��-�l{�xy0�.{yם ��w���Y��# N��ɽ�*<eɽ�*<eɽ�*<e��*���FC���;8�jɊvx�4�b�z�a�"s1
�5�Ҟ\�ռj�|X���Rr�ӕ���cJ}���޵7��j�Р��%�u�){K_5�M�;)��A���S�Ƃ��ɽ�*<e��*�������Voցt+�5%�V�²z<rF��������B֊ ��f��2�a�D��3�Գ������q�j(�d�A��S�Ƃ���W�'�㵥��}?��D�����G�k`>-:E%��D�&t�ؠ0v3> � 	��#�uX�����:@�y�v�Zɽ�*<e����T�����W�u5L���j�Р��%�u�){KVMr2�����MS�������
+C�˾�� ��*��t Եp��r^�QW���B֊ ��f��2�a�D
��
���t�U�Y "�t��{d�.{KP�^�%� �F�_��Zg�a�J���J����j�Р��%�u�){K�G`�,�CFG�؍N�qGw9�Yzɽ�*<e��*��d���=,�o,�����5��[1gSD+�?M�וۏ�¾-L��vYw-h�(�Iɽ�*<er���4GH�)^۞�;��޶(:�B֊ ��f��2�a�D
��
���/}�	�S��ɽ�*<eɽ�*<e� �F�,$�`i,0����2}x���Q�px����Hk�K{�Ե��������8�z�qs�ɽ�*<eB�/k�R1RMQ¥���`�k�hE�����V7�@3�w�K�Yc��� Nb '�8�)&�0_l�u�I%�F��A��@V=����2}x���Q�px����%���NbqB��z'OΔ��B���uFS��4��!1V��+bZ���1�0�.{yם ��w���-���Ծ��� ����~�XkT�0�� ����~���M�Ϟ�(c+~��ͮ{T_���ju�b����B֊ ��f��2�a�D�ި}E](����Ðjs��Q�zO�;8W�f]�bܲ!f��|835� g�4�u� ���5��[1gSD+�?M�cM堧땂�C �7�
-�yz��FS�Z�:����$aځ����L�����`�k�hE������5`��d7��VZ uD�'*F�l��ɽ�*<el�u�I%�F���[Le�2��"��N�v��,���A)�^U��R����+�6t�m�Mc(J ���I@T�ތV��P�����|�kG��[]\c�mؓl�fD�1�Jn����4�u� ��͐�������O]\#����r�}�S�axV�\����i�}��+M��?I����� 5��J���lZ����\#����r�\ `L���PY4O�L{IJ��n�Y9⓷F���t��xl�	!	�6��䀘�4x}���Q��^5:%�||lu�P,�:S��]��-��H�T�i���t�4��()zӺ_gR�6W�mQ���=��"o��{�s4υ�-J�����l��,���ҿ%����D�
2��C0M`�%�hP��d=MK(�b�sN��8H��ޛfe�^C�ɽ�*<e�����Q�`~������O��:�g�'��(QC'�K��w��G`�,o���R�-��7k��J7�����K�am@�p���b�!����h3���*�Ӈ�k���,(nɽ�*<e�VR֒�;�Y��##0��W�d���C�^a����Rb`x4����p��ɽ�*<ev�7�w��t���If���9TI'�09k� �f{����2#_w����]�0��\����i�}��+M�l� ��&��5�MP��px����`q��Z�7U�'R�ɽ�*<e �.�Qq�*����p��ɽ�*<ev�7�w�n��=)�'ѥ䰾M^� b��pXd�4���Ai�"&#�����n��;��2��:7'$��R��e�����kV��q�И�mJ��E|�m;ɽ�*<e�����Q�`~������O��:�g���L�d�_xZ��C��5��I�A���[��Ƹx���]L�Eɽ�*<em�x�˝��i�P�����f���9TI'�09k� ͸!Xa����dGUĖeU�}x���Q��+�(�T	�ɽ�*<e1��0����,�4����0b��*��-`������F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)X$�j���
&��.����b�g�V�����F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)Xh�>�(Q^9z(r�Q�)RZ�]�,\(�%d9�Oe���<]ΐ�i�+��j�;7_^�LK�ŷ����X��X��O�
����KvB�"��A���=��Z���ZT��6���w4��k��O107���z��Y�����p���z3��R�wY�%Ls���������޶(:��6^��a����kN�~33��_���S�픺]'E���iu��Ը����$K�
��ցt+�5%Ta�upI�]'E���i���~�U�j�[<�0��\#����r��4�b�z�aj`▘9Ё�Y�`��>�M��)����n��d��)%��b0��a/v�sݏ����p����}Gδ�-��$Q����x���]L�Eɽ�*<e@9_@�R4�8ߜ�R��ڇ
�܎[�H
E#LPA�Y��g��8t����Yr5�_F��x���f�2�&@y��Ų�.����e����NxL �?ȯ�r{�Þ�{r���p��$K�
��ցt+�5%�ʬ.gx-�P���Ξ볯`A��ɽ�*<e��}Gδ�-�5�MP���^tD����U�y��7%Y�g�E�#������Xƻ�2��H���I~"ʒ�������C'�K��w��G`�,o���R�-�_v��G�]��/�žCɽ�*<e����tW���O]\#����r�{E�6��h#A�Y��gɽ�*<e3ƹq�nNs�/��Z �^���<���^��c��d6ɽ�*<eɽ�*<eƍ����3}��+M�C��\@���
:��{gɽ�*<eP�7ٝGy�ɽ�*<ef�{��t�'$��R��e�_o��u�����h3��s%����3JПE�[5ɽ�*<e��E�5���������V��F���2#_w���r��j��9I�3���ytp�^(]e����j�M��Eo�$g��ϫ���~�Q��u���Yݿ� X���K�ѥ䰾M^��i����1y��V�7UvS+ё@a����kN�~33��_��_��q�wY�%Ls�������J�4r�Y��X�Bh�W�	�y{I�7q��]-�s�eS�z��z\#����r����#h���h�q��$K�
��ցt+�5%���X�u÷t�4��&*�w'�-��y�s8�SV���y���՘H��	�e�]�$K�
��ȋ8+�������p��́�g�N��k��O107�% >��^Ue/�G�U_��YE�g�%�b��&��d��.l����r�g/�G�U_U(��T�u-�ɡ����������-�V��Nu:׈S�yg��VD�j`▘9Ё�Y�`��>�M��)�atBҷ��c A�[f�矑��ӆ�澮/�žC��
���UcjoAh�q��m!�qɽ�*<e���h�q��$K�
��ڇ
�܎[���҆��A�Y��g��8t������p�� �.�Qq�*�`V�f�Bɽ�*<eO�
�����ASJW8Ǿ,GLY/]�������7Ց�X2��~`��r���-�rS��8��A��(Ѷ��$B]Qx���]L�Eɽ�*<e���h�q��$K�
��ڇ
�܎[i�j[�r��;7_^�L�s�C#e�uɽ�*<e����,�4ɽ�*<e�+�r��y���8t���^�%���ѝ�L��Ԝ�#|���;�ցt+�5%��J`-$�*Χd'1�r,\�����e'4M���/v`S^!�������f>>_YRcy�P����*D!ϝ���g�H������3\\<:��6I �I��ѥ䰾M^���F���oI���ܔ2��t��1l��Fx��ʡ���_��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e=��d��p�^(]e����j�M���;eXv>����p��́�g�N��k��O107�% >��^Ue/�G�U_T���N�LZɽ�*<e1��0�+�r��y�Q���'�}�ٔ^qt��DzjڢXeS�z��z\#����r�LL�6ۨ�V���F���=Si�.��ԷGс�	����сZ4�Q*#9?��{�h?�EG�1�p;�@��6�Jx���C�U�5�MP��px����%���NbqB��z'OΔ��B���x;U/��*�����Zɽ�*<evS+ё@v����t\Y��پ�?w����Ot�;�Y��##0��W�d��y�ֶÙ)ٔ:�OFDG�@<O�G3��6���m�ჭ�u�l�d��WX��P
+^��OL� l%n[8�q��Ӷ�;�Y��##��F�<���4�d���s��Q�zO𕓔��m���	��V��P�����|�kG���p��;��U���W��)�8ĺv���-��i� $�cr�j���%�a�9|��ި}E](�h�#��IJ<���	��+W�L��W/�p.�qG�k`>-:<�������iP��[Pv���-��i� $�øxQ@Q�;K�N��u��7-��]��f�|��R�OO���T��<�n�\\#����r�T��w��7;Ĕ���Í�ǕvEGL"~_D��D�i�`"u�y���m�B����L��()`S(�K{�����Y�_;���%�Lف4c�>X�������_�<��N�d�)f��X����"U�8?1A��!�(I�Ԕ5CIE��LL�6ۨ�V���F���
��
���
EÎe?����mv�ۯ��1�s��<��G���"���}�Z�z�z�LALƒE�I6��mq�\F�Q$=�u��Z���1�����с��֎���\��}:�f���L� l%n['�=�3���z�%̗��mq�\F�z�a�{�s��
��R'����сɽ�*<eɽ�*<e�C�\h~�5�p��iZ��J���J��RKD�vQFɽ�*<eɽ�*<eƓ�pp��N�,�|[��ƅ�������F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)X���9��%�EX��Yj�>����z��]�Q:S��]���v:��l�ŘP%��ޘ
���FB8����{I�l�UY��	r¬���{�#�C[+,���tn�~����i�}N6�9_�[��f�c̟1���Ɋ�|��p�l��U��h�\H���jdqko:S��]��rX����ȫ�$m4��ji���q���Y�r93z፥ӕ?"������A"�1֦��IPs*�:S��]��nfph��T[�'2:AR���=��a��o��<�gf3[��;�	�-���30�\�0�&�7O"�B��b>/��2��TȞed"��d������C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S��(�[�v��6��D�SG����jp]� yR���g�M�9�mćX�V�?`�I=(MX�*ɽ�*<eɽ�*<eɽ�*<e�C��ֳw�^;�\��^�s�H*t�ؠ0v3>#"܇a���DF��L*+e8`�q}��+M��gA�=���*�M���-���Ծ��#��V��9�=�G��Yr5ɽ�*<eɽ�*<e�ub����T�2+��@�l�VUQ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8������MP��J��3��HY ����3\�!ќ΀y�U�I^�*^pc�cJ�� �4$[��)v����Ah˒�1:S��]��/��Fs'���\����6�����6)�$ˤߚ�(^�^ ~�I1gn�m^.��?TԽ0�1���Ɋ1�PST2'��ևc\��FHx-��ƎH��8�盕k�[��C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S��(�[�v��ǯ�� ��7Ց�X2�ѥ����xE�p?��7Ց�X2��~`��r��ײz�'����jp]<7� [��ASJW8Ǿ,GLY/Xƻ�2��H���I~"ʿ�,>)��H�"Uy��\=�B��YXHv@�������!�f8��aI0��GȋMFx��"��DzY|�;䋄C0
��Ɠɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��*����*�M���w۷�Γ��K[�k�&�r���4�b�z�a�"s1
�5�Ҟ\�ռjW������%�F�h ^'Ŏ��Gb;�V>�Vt�ؠ0v3>�˯.��s��P�C�eD�8n�ɽ�*<eɽ�*<e��t�F�f���9TI�;�Y��##�1{bhA*}|��rA�Y��g�t�R���@n٣�r��QӚ�E��dd`�(�M:S��]���3GI++�ub���-���Ծ��#��V�;0c���]:ɽ�*<eɽ�*<eɽ�*<e�Be�����C'�K��w��G`�,�CFG�؍NI�R��
���V>�Vt�ؠ0v3>#"܇a��[�r��H�ɽ�*<eɽ�*<eɽ�*<e8�q��Ӷ�;�Y��##0��W�d���C�^a���w�E
��Ɠ!m+�V��v�`rv9��A��/M����bɽ�*<e��*����*�M���-���Ծ�`�� �P1s�1��';U�`�� �P1sRI�c�@�V>�Vt�ؠ0v3>�$(�dOYD��ˣ��Ez`r��ɽ�*<eɽ�*<e8�q��Ӷ�;�Y��##!m+�V�e������e�>��9�����Ym�z�a�{�spx�����m����k]����5�#e+�^�Liɽ�*<eɽ�*<e9����`�n �u�HY
�H�8����{6;IFRq���cQ��y	�X��ub���-���Ծ����.ޛ��.��O�����tgv
И����ɽ�*<e�Be�����C'�K��w��
Oo��"/S�Z�:��]j�=d����~�1�7
�X��d,4���?wn}y$���:�g��7-����u2˙�-?ہރ�ub���-���Ծ�6�_� �n�ϘV�q�e|β�,Lx�ɽ�*<eɽ�*<e�G�OLJ���
���2A�Y��gi��k,��ި}E](��H��J��ި}E](�M��hBM;ɽ�*<er���4GH$
?�؁ޅ����)iy�V>�Vt�ؠ0v3>Δ��B���]4�vj��=�E�I6�'*F�l��ɽ�*<e����{����������UY�s.�|��,���וۏ�.�E>2�<U�S�Ƃ��ɽ�*<eɽ�*<eɽ�*<ev���-��i� $�\�`�P�J�@.��X��d��*�M���-���Ծ��#��V�C�2w��Z[߷�J��A�Y��gi��k,�
��
���t�U�Y "�t��{d�.{KP�^�%ɽ�*<er���4GHc��Af�̠o����4�b�z�a
��Ɠ`��ζ?��Q8�斆P��S�5tV��^���>�A*���s�HB:S��]�亶���ΘA�Y��gi��k,��ި}E](����Ðjs��Q�zO�;8W�f'*F�l��r���4GH�R���&�!�^�BOP�p<�G ,4���?wJ^f^�A+�[�	ݛ� ���������mZ�ä�A1���5.�8��?�RY�z�a�{�spx������JFV-O�;8W�fn�������rt��l�-�B�N���9����`�n �u�HY���W�2�rt��l�-/&6C_��SuJg��/.�w <>k����$�ܠ	���Ɔ��"�����F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)X���FS��)��|]�zg\�[Ak�mؓl�fD�۹:��'�����5{����vA�P�ɾXe�g�:4�Ee0�q_}�Y�[مi�����>�m/*,:�^�5�{�Ѩ����2 i�ZO�)?6����L<ިq�>��1H����T��᫞e-��1�~��:�@i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q�݀Vh��5��3}��d��p�dGUĖeU�b��i���sX!�_Өg%��>��fg6	xɽ�*<e�/���%�N�@�>=3t�끆E�n�P��Ti?���6�:������ჭ�u�l��&��>�^j�w���#�%���ɽ�*<eFª$�cJ/���<�������y�|3k.sb}ɽ�*<e]�q���~��_ ��끆E�n�����Q��F�g�pζ���������s���4T������R���zg#��AD8��d}���DhY��F�ɽ�*<eջY@f����cW�Kg��@հɽ�*<e"�Y�n����3WWC�5�R(�*��؊��SV8��+ Z��L�B"�MlZp
T�m�B�������Ec�끆E�n�r�=_V8��+ Z����w�ՠJ7�����K�am@�G���L�w��9��V�n..+`��ɽ�*<e�ASJW8Ǿ,GLY/]�������7Ց�X2��~`��r a�����O��:�g��K,��W5�R(�*�������ɽ�*<e��L�B"��I>/�4	B��@ȏӽ��9��V�nŨm{�2`.ɽ�*<e�ASJW8e����"Rݗ]T��~a�2�]ߪE�g��EڤoUx�$_'u��U���mǹL���A�끆E�nC�Ѝ��7]!�{������w��7�pI�3*'K��>.ZU�끆E�n�)�	5G����՝���џ���2TQ�U7x"̠o������V�uCM�Q&�"��q�|�"�����/���%�5�MP���J&K6���
�ޘ9�v��̟�}3��|��V8��+ Z3i��b��̸B�����{���̙�v��̟�}����%�#��U��Zo$Ԏ !�\V8��+ Z���V�uCM����C=����P��/���%��R����+�6t�m�Mc(J ����+�Cp6�N>��Ӝ�TO�Ɩ�tzɽ�*<e��]�Ͻ`�N�,�|['�݋	��`��%-�T���}e�ɽ�*<e�(͋�xF����v�7)�"Rݗ]T��R�W��3N�܇���`��1N{� ��{T_���j��d� �}�N>��Ӝ�� ���+�'V����;� ��r	(B&0����cW�Y9�SGiWw�҃b�a��b�y������t,"w���[7���cW�Y9�SGiWw�J&K6�	�밮�:�g��7-0H�<Oa�B�_}ʘ��U�H���jps� �<!F2]�J8�F2]�J8�F2]�J8�F2]�J8������MP�_����be�A�����;18�^��F��Pj :S��]���>s~S���i���8�(KpJRR��蠍Q3V ��zU`��X�6ƌ�f8�:��l�щ���-(?M7yWPI	X���J���B/�E�d:S��]��Ù
I8��\��د8J�$�
)�/<�����gֱ���\�UF2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^���9_ߏƮ�@���[��ў�ѶG�0���ZEM�ɍ|>�G��*�20������d�*C_����,�g���U˭4p��~~�Tfg.{��f�r�"�: {�q��I��/eA�k���	�F����9���rzM=�z�j"��w8Oy\}��:;����{�/�d���(�-����)P�hx����ʢ���f>;�݃����h��D�O�������Ù����6�cW�n2dꜱ+�	hp��Ԁ�F�Y���~N��g[��B�s(�?A�Ҏ&�Ё?m�-�,�X�Ÿ�f�2_B@�~%.DI���:��t�%2�/	J��hא�܇*9�2�\c�5��u|R���GX��a��Xڟ3�8�H�d�h���� I���}�t�wI'[]
*�J���oE����:��C�$k5p!,�7ڐ9� ��h��'i沃�Z}����Hc�9�%�\T|Aů� �B�#��t�(a�����z}�E!Ͽ���!Lؒ&�bL�.��. ����lB��,zyj���0_��A�\��B�N��%졖*��j)?��(a�����@��$�G#�ӵI�0��#Ҟ�s�-I@>������BP�\_�0'���I"ʈ�W�rB�������i0aXK��2��H����D���i�6 ��Z�)a��\ `L���c��}W�R�#C,��n�Yx���|��/_��P��r�k���g��� H]K�s��K���{T��
�7`�	�6�#'	��m�:��eH��J�	��[W�DC�"�N�?�ot�'��#~D��\��KB����VL��'�s���7K�f*���b�0qK�s��D�1d�	!4wI�o P��z9����D�����e�mu���H��H�
:��p��؋9i�^��,1DԾ����\J���H�.'a:�s�c�A �Ы���VI#�1z���x�q��Ǝ�b\[��½�#��$̆���5��0^v�'-�r�D��6�^i~��b!�t�&��9W����m�$��m�?�0.܍�G.I�TVzi C�"4D�MUP\�0W�1�5<�蔺Z�ØKϔ������!1���s�D|�����N���Q�)y����:6ݑ��/�^�L�Lr)��ש0��b=��K�X��u�Md�����g5m\5 �Β����ܔ������^u�{�=.��x�bW� ��:���ƺ#�FE��7�R�b=�D2�F2]�J8�F2]�J8�F2]�J8�F2]�J8��ې���������U�F�/��f��i��˳���}�]�v����phl_>וL_g!����8�'�-�pE�.�"�$�'��!�i�uc�����F2]�J8�F2]�J8�F2]�J8�F2]�J8��A�2c�����O�:���<��	��^L��C�;��,�7C	��ṥ �u�o�o��|��ʽ�|~%�������&�U��uSF��~�G��1�)JO���ĸ3���ꤢ˸S��ƀԫ��	��ߟ��1(K4��.�� �|�D��!���O�������Ja�]_�A����n6�8u
���+��֮)۶�4����E�����Ǥ:�P�%U�Qׅrڑ ��-���@�f�7zX0�k��ܷ��W"Цe�?�PX�Z��J�;=�d���{(�rZ�������F��܀�TF��%��H�E\�J����L�1��8��Ȱ=�=[Ak�N� Gm�07S�&A��Q3��w!A�֌�g:�Bح������A	s���B�p��3Ԅ���.�?g��3nQ�XzP���`j�{=�}\��8B`}��t�q����DF��t37�h|MH�����z�&��E���ޘ ~��fɽ�*<e�N{}���m:~���J�^*���ɽ�*<e�N{}����'Z�Qln�5Ǔ��G�tx�E�Bx ��J�e7��e���>sK�EbcW����]iL�<�@T� ��t�78sK�EbcW����]iLVB��*�exctw?�:�=��=ʱ_p���X*��ڳ�/��I�U�Z멿�*[���d�n��Q�DjL�b�Ff|Iz�c����1S��M	�I�.Q"-Hw^��蔂p���{��%W���h�J%�Y��Hw^���'N	�֜��%W���h�J%�Y��Hw^����uۨ�T�s�g��8Z	�I�.Q"-��X{m����rZD�Q
lR��RT�Jl�4��wy f��F=mOu�r}�I�tsC�0�~����~�M+DW��-mL�o��1��UC
��ɽ�*<e�M+DW��mOu�r}2�֑]>��mI�z�#-K{*o��^��tL�
����=��Z���s��[b���x#�"�U��xRQ��L a*�ĭ\Pһ�I=��R5�+ұ�i�A[�%ѯ��a΋O����E�们e�c]���s�c�����"-w��-�'Z�Qln�5Ǔ��G|3k.sb}"-w��- ��01�7g �9bA��ɽ�*<e�m���g�q�?D��\�MP[7��͸�R5�+ұ��d�':	�{��rm�����5�3P�e�[�[+ɽ�*<e����X>~A�Z�\�|���L�N�����]iL��A�|a��V�)�qJ�^*���ɽ�*<e�N{}����8�����t,x�Ik-��.�ֱ�r*�M�D��~^-Ct��Q^U>a=���ھ��:^��ġ��N���r���4GHvS�축e.M$-����BX��hP�A~�$r�0�2���*@:�mc�oK�~�E�~`zR����KDYn���{��B/Pb��|�\��7��r���4GH��^+���f����u�J�[�[�d���7�y��|�#6�=E�y�m4�y�����F2]�J8�~�&T�S�۵����0��m��yQ����Ci�ܛ�|�F2]�J8�	C7��3�^�X��]��zN�����ɽ�*<eɽ�*<eɽ�*<eT#@�GN&I��rU�Z������ɽ�*<eɽ�*<evS+ё@��n��EC��ଡ଼�F2]�J8�F2]�J8��C2=iO)3����phl_>וL���ה9������F2]�J8�~�&T�S��a->�d�W�����D��5�3s`�J+�ag��*Kv�����~.O�~�e�U�yl2�����C�g�V�uۨ�T��,����n���)-:E�%_1W��X�����a->�d��x��{ɽ�*<eɽ�*<eɽ�*<e�-�YR�)squ�`�)�X��]��zN�����ɽ�*<eɽ�*<eɽ�*<efMT�Ҁ��H�ڸ��P���S���)�ߴ��BYA���L�N����,����nd�sߵ�=~�[�eonD[��]��{(W'4�l��u�
�l]:G�&C���~��ĺ����ىn������J������\�X��]��zN�����ɽ�*<eɽ�*<eɽ�*<e&6��u48H�ڸ��P���S���)�ɽ�*<eɽ�*<eɽ�*<e!�4@�+ɕ?kV7�(��^o�&I��rU�Z������ɽ�*<eɽ�*<e���F+�N��S����*\@n��{���}Hj�w��p�@�ɽ�*<eɽ�*<e%ߒ#@Nܿ�P�6;7}q�cW����5��M����|��mHɽ�*<eɽ�*<eɽ�*<e�c����Ϛ�9����	��y����}Hj��\�S����#�Ε�@�>֠�%ߒ#@Nܿ�P�6;7}u����v���}HjIe&�A@ɽ�*<eɽ�*<e%ߒ#@N��������A���d��X��]��zN�����ɽ�*<eɽ�*<eɽ�*<e�ܚ���ԯ�f�y�����Ќ����
�a���UUJ ,�z����e+ɽ�*<eɽ�*<e!�4@�+���(�-����)P�hx�d{.�D~��5����fF2]�J8�$�䠢O)XimϿ�wz�/��Q��ѕ���sg�vA��R*�D��|F2]�J8�F2]�J8�[��ҵ�UUJ ,���jcO|j��ޘ ~��f&�r��VU�	(�� �~�e�U�5��M����|��mH��z: �7��<���J&��Y��`��;@�M6M��1���͛5��M����|��mHɽ�*<eɽ�*<eɽ�*<e��;@�M6�紻�p�#�]
�����e%�ɽ�*<eɽ�*<eMͿ���q�r���-���W<:K@�[G-sڸ�OB���c��LL�c&�r���lև4[@.Qu2T!�қ5��M����|��mH!���dT�4V{1E�I����=�HP�N��||�,�h{�Zr%����g�� }�T�����]v��sK�EbcW���,����n�m�$Τ@��n�W�DA_:����W<:K��S��Cɽ�*<eɽ�*<eɽ�*<e-ʞ&��J�c��<���p�"��f�:.H.�4&ꬶ�Rɽ�*<eɽ�*<e{��<Ia���_�av"O���#�]
�����e%�ɽ�*<eɽ�*<eMͿ���q�A������s �� o֙n,(�H�y��8d�%���ɽ�*<eɽ�*<ekwO�&뿃,�M����5��M�����x��{ɽ�*<eɽ�*<eɽ�*<e���3A�^x�ɶ@�F� z_.?�PZ������ɽ�*<eɽ�*<eMͿ���q������h�^�K4���֢���N�������Zɽ�*<eɽ�*<eɽ�*<e��ǔ�7�_�V&IM�f��QM�g�� }�T���a�;^<q���_Y7�{b��D�:�]�,VD���1�k��a->�d�|��mHɽ�*<eɽ�*<eɽ�*<eך^!NH7��z�IYLy���k�L��'XD?jy8�e%�ɽ�*<eɽ�*<ekwO�&뿃�jHi��^�䛓��yl2���@�[G-s���?�M�ɽ�*<eɽ�*<eԃ:iD��z����ت4/�s��"�w�UUJ ,�z����e+ɽ�*<eɽ�*<eY_���7��M��c��xÅ���(�xt��:[&I��rU�Z������ɽ�*<eɽ�*<ekwO�&뿃f@��S�c��.�$� 8�(��Y8��W`~��Z���/^���$�ul&�2������N���[v�yl2���;�e(<�KB�hE4�`sm� 7maH���	3Y��
���|H�Pk���,(n�����I��嶡+U�n)ɽ�*<eNM�\�*~��?D��\��.����iʆ�S��3bc��?�C� e��ejр��?�C� eY��$Y�aھi��͗
�z���^BQ�D�o؞A�Y��g3��֪���X���6�\��D���C>��M �IꜦՕ�P�pp-�͋��#��rW�0N�<�|a�~a��SW,�̼[i''
��I�q�D�&�|�D������O�g�k��%��&�|�D������O���x�&:���
����`r��κz_��d��t�����Z�\Ȣ�D �.�Qq�*����p�� ��� ���:�f
�{��t��۠�F���:��nB�r�rz��Ff|Iz�c�jaq��݉#^ͱؕ�͔����Y���mf��uВ����E�
k�m�Ϥ�<y?��Z&�mW���JYw�8�r�rz����p���{�C�e
����'�S������Y���mf��uВ����E�9�Gdo�03���р�"c���Y��@�đ�k��S�#���,0+o���7!^�߸�'�S��!����f)�e�>��i�f�j� ku-� M"�:�KD���RI��;�!1�0BۀZݪ+i0�6B������"Rڻ�~P�� _��?-�)f�T���yTظÂq�Ff|Iz�c�jaq��݉#��9�4�!X�=h1TظÂq��uۨ�T紊�y+6��9�4�7�����?Zݪ+i����������
�9��%������W�����;�X���A���qvjV���"x����lafG���k��S�1O������F���Y���^�֦J��9J�W�U��
�؃��Pͬe�c]���o^8�2��弯���l�Hi�X&�Mo�H!�|�G�S�#���kp�P�)��\�u��y7ɽ�*<e}ʈ \�/He'%��@�|���ɗdW�Ј�Q�7�c�Z��U!(&>,���x����u�~zbF�j�����p��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��E���ޘ ~��f�B迸Ψ�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eQ���v�&yu")�
B�pe��*qb����J�n��e�3��:uG��u6�Zݪ+i���������Y�R�GL	��D2L(��T}���}�ʳk����V��+�
h¾n�5Ǔ��G+o_�o������L�N����l� ��7�d�'��O����ɽ�*<eɽ�*<eɽ�*<eɽ�*<eڨM!Q��s�m]��ȋ(Plkɠɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�Z�\�|���L�N�����OUi�_Zf3�����^�֦J�����a[�&x\��斳pچ��zsK�EbcW�yu")�
B�_���QR�{���lU�W�ee�u����Z����sK�EbcW�a�����F�K���آ� m���kA�Z�*M�RT�'d����k_�j#�.��zY��`�J%�+ŮMW����/�K9��gCf��¦*��dQ1y]��%��D�d܁�v�lˣӸ�X�p�_����n(L������7FC��_�����%��0��P�줆�׻;��O�t�� Y� m���k�F���_�|3k.sb}Hi�X&�MMj��*2j�n�5Ǔ��G�W�X�u{U�~L�?��{v��ᄎ}�ʳk����V��+w�u��V|"�_엘������_��7�>����kN:>և�d2l�}�ʳk����V��+gxZU��f�C}�/��cV���5v3UF2]�J8�F2]�J8�F2]�J8������MP��%�0=}�����I�T�ﭦO��,���V�i�s&�*>ǚF2]�J8�F2]�J8�F2]�J8�F2]�J8�*����n4Ck���nK����l����7\�~s-����ԙ�7�b�n�;�o$��q�Qy[�^N{�<�R�Lj}���t˥SH�������h�fd�	m�L���W���F2]�J8�F2]�J8������MP�m����>�ɡ3@����C��nhV���5v3UF2]�J8��&Ic�E�J*RK��s�T�=u��\\#����r�׌��u��Z���/J�!#�]0;�G�	�M��)����n��d��)%��b0��a/v�sݏ��Ę�c�����N�ޛfe�^C�ɽ�*<e����m��b ���@��l�:iF]�x����cT��%zؕ��g�q\��/�žC:�]�,VD�ցt+�5%�D�%uޫ˩*��%��T���N�LZu:׈S�y�է '���z�6|"��K	~�������4w��������fuh�+�fKˍʔ��j��ej���/iԣ�֎%;���['$7��/�žC!�4@�+\#����r��y��ej���8t��}�tؤ�l�k���,(nO�
����'�7� �EH�S����{����,�|&2}��$R�������٣wc����p��%ߒ#@N��������G'����ȋ8+�������p��r�֏��9��W8 �+N�����p��%ߒ#@N��������G'����ցt+�5%�!�/vx�����p������,�4P�7ٝGy�f�{��t�b/d2��s��f����M��c��xÅ������`��f@��S�2KG�E���j���(�[�v��Ls!�EŬNl�>*�2�G���_D`Ȩ���QrNl�>*�2�G���_D}�S�axVF2]�J8�F2]�J8�F2]�J8����"F�^|��]`�O`��a�R����>W�_����N4�F2]�J8�F2]�J8����T%�g'j`▘9���~
�l������V�3yn�3���IE�گ��L�����Ȫ}�0)��bhF_8(uR�|g��b\	y`�!���dT�4V{1E�I���䞈E[� ϫAu���T����W&�x���]L�E��9�Y�X�B�$D./�j�Y_���7^|��]`�ي�L�<T^|��]`쮤z: �7��<���J&Q��>M�<9�ݞR��=ӂ�ѱ~C�F2]�J8�~�&T�S�W1����1g��M�b���S�/�����C��nhV���5v3UF2]�J8��&Ic�E�@�[G-s��5�3s`�J+�a�a`7�v���\˪�����
���2�=r��֯������śt�^���� ��}���AEٜ+������ވlY��"D̢Д�٪,a��(�ݦ^�yl2����s�]o�<�<�Z�%�<���J&���y�<xu�[0���ߔG�=��y-�JV;D:���Ŭ�+�g���śt�^��Ü<�Z9�o]н�������r���c�K��b\	y`�w�fRԾޛfe�^C�ɽ�*<e��<RK�r�M)YTs'$��R��e�����kV����Ɔ��"��<RK�\�w�:�	��FLE+����kp�l5�*N�sڸ�OB���c��LL�c&�r��L�#�W�E<��	� ��v��������?�ɬP�e�[�[+E�I�����P{v?�f:5�5ǩ��'4M���/�V�W�v#@�|�0�']_�@[��]�|tֿk���,(n�|�2<sq�l�Z)^��_�����¡~�x���A�X���(����F@�����p��:��8싄F�p��#����tU��u:׈S�y��L��Ԝ�x���]L�E ^���F۴�˾�[(Y�2��a��[�eonD���t=�)ɽ�*<e�p��S	�ȹm���6�"�B�b�[��7ɽ�*<eR}��G�<u��rnN�-����p������p���P�g�c����&:�A`�l��e�8���ֳ���$]s�m]��ȋ�#��VХ�l�/޽�'n�5Ǔ��G�شM�ў�NfMܖ;d7
�n ����
�9��%����e��IB+�!ɽ�*<e���7	��l78����٦��� dF�R?��(�v>���yu")�
B�K�]=��"ٰC�QS{Ԃ9Sfֳ�-�V���ZMD�
�Ύ�F����J�n��e�3��:��5+`I�'$��R��e�����kV��+�r��y�9�ݞR��=��!5��tl]:G�&C�mR*�5:�G��RO��ŊN�:Ll�{;Dj`▘9���~
�l�������G�?fT�ܹ��J�o+���"�H� ˯nkB�Js�eR��_�`V�f�Bɽ�*<ey{���V5�����&q!k4��3��^&�|�/*������J�$��D9� 1ɽ�*<e��\˪�����
���2�Pn�M����
���2�UV�ː�	�*\ɹ����LФ��sK�EbcW�yu")�
B��a[�e.y{���V5S�%cd:�io�^�ơE�Q5����X��0h����8t��}�tؤ�l�k���,(n.\��O�dF�R?��(��7O��L\�� D�4I�FQK��v��,��MͿ���q���
���2|��chRL\�� D�
�d5A�3���UJK�R�e9k�Q�yu")�
B���l� ��;Iyfs�kp�P�)��شM�ў�NfMܖ;d�w�Ey�@��$l��,\Pش��M{a����x�^6��u���S���,\Pش��M{a����x�^6�ý)����A<u��rnN�-��+�X�{�{��<Ia��w��\����)tK�:5�5ǩ��
�9����'4M���/=�B��YX*3ZC�q����,(Q'ƃ�l��C	���D�\å�o��[���ޚ"\��ںy�#�)34*�� ���
�9��%�����B�.'7un�5Ǔ��G�شM�ў�NfMܖ;d�w�Ey�@��$l��,\Pش��M{a����x�^6��u���S���,\Pش��M{a����x�^6�ý)����A<u��rnN�-��+�X�{�{��<Ia���[�eonD�+)��n��c����&v��t�c�9�ݞR��=�ֈ2t����`V�f�B{��<Ia��?)��O��6�S��t0.d�չ�R�l�VUQ�F2]�J8�F2]�J8�HE��޻'&:#��M����b\	y`�@ػ ��*ۄ�y�	c�i�ܛ�|�F2]�J8�	C7��3�^������Ą�#��MͿ���qzGך/���b\	y`�B��OS��UP�h~��L���@l� q����d�v ��j6<������J�=aS��śt�^ۧ4�a�ڔ�~����҂
�9����C��ଡ଼�F2]�J8�F2]�J8���9ަbq<M�L>�;>c�ݒ��5�.���7������F2]�J8�~�&T�S��v����ZQ�R�"=�{/��f���D�h�*���m��Lݴ�����ȉ=���g�H,$�`i,0�+j�Lp�jHi��VL�����]T,�����nX���Pbg[����9������^�M�/,�mV�*���m��`�C4�����4�Z�
�Gc�Y|�0�÷���������F�Jz�j����~�q%�e�T	��<��ͺ��_~��]�)�{��s�����ߪ���
6ţ��|���P1޸�7ka�`eI��/�žCa2�C�8�W�a/v�sݏ����p��;����˯�J�(q��NIL�./�j�"7�!ne*5M�L>�;>c���.˟\,�Ҭ3�Ss���C
�V[��q�И�mJ��E|�m;ɽ�*<e�=��>[�{��y�a��L�T�	�>�D���7�W�Y+� �#
},M��j��˪bc:�^�6C_ZWA�Y��gOj��cI}3\��М}��(H��u�6����e�>{И��Cni�'\�g�i�����7vɽ�*<e�R���b8V������8���L�8j�!Yn��R�ɽ�*<e�S�Ї1�lr~�F��[˷�*��,����تa�ɽ�*<e���L��nj;T�:Nw��Ҩq����H����nj;T�:Nw��Ҩ*���qT`�&Nꊓ�Hb�Tw��� �^S�n�Ir=Xl��.苢��w�MͿ���q��^�e"�r~�F��[˹�`�7.\�Y�=�5G����D.���nX���{��<Ia���rq��&��B��)���Al�'0�r���4GH��o�ȳ�Y_���7M�L>�;>cץ�|(i���Ina�_��M{/�� E�^��U$/V�b����9��t�|J�I�?7���_��Fn�p�-W4+HS�&2�y�*�h{�2���e�I�v$3|m��X4:Û��ɽ�*<eLݴ�����ȉ=���g�H�˅&��E���
����M��Hn���X���2��5�"���,}v�͹j���,�.s&^�mJ<k���,(n{��<Ia��<X�3Ѧ���0})dT@�q��+�Z��!	�Y��'N	�֜��%W���h[��x+�fMT�Ҁ��A�Y��g��9�Y�X�ͥ�1>���j��˪bc:��ae�ʳ��s
zl���K�p��bxA�(N=��B{�]kKE�����m�6Ī�����8���L�8j�d�������uĥN�$L�_��D1A�Y��g/V�b����9��t�|J�I�?��bV�Ƃ�Ԧ�0}Ъ�����8���L�8jr����Q�:h\rһ�����gZ�M����p���(_qn8�P <�t-*�*�N0�<T��*r��|��Ԧ�0}Ъ�����8���L�8j��qz��m�U��GBM���gZ�M�ߔG�=���HQ��~�,( 9������p��{��<Ia���rq��&��B��)��$���{�8�ZQ�R�"=�{/��f���D�h� ��㼽|lɽ�*<ezu�V����ɽ�*<e�(_qn8�P <�t-*�*�N0�<���m+�%`��rq��&��B��)���&�p�2=�*�1��v��,����
���b��4ڠ8��UC
��ޛfe�^C�ɽ�*<e�X._�� <�t-*��HA5CE���9��p���b�!׋q�И�mJ��E|�m;ɽ�*<e�X._�� <�t-*��HA5CE���9��t�|J�I�?��&-�ɚ�9������^�M�/,�mV�A�Y��g9�ݞR��=9�ݞR��=�5����fF2]�J8������MP��{�'͢�@ػ ��*ۄ�y�	c�i�ܛ�|�F2]�J8���e�̣A�̌N֓���~��K[�k���Tea�T�=u��\/���?������ҥя'4M���/�V�W�v#@�|�0�']_�@[��]�|tֿk���,(n�|�2<sq���c��d6{��<Ia��/���?��c�����Jt���y�PAN$(��5ɽ�*<erj��`�^��h����5$�`o*���N�`?=0.d�չ�R�s8���1�"�ȹ���/�žCr~�F��[��O���}U��P�8�z�4�)11y��V�7U^(�v����$r�0�2V�NǺ���-#�6f ��V.�˸�k�7�ղޛfe�^C�ɽ�*<er~�F��[ˎ�Zg~���_M���5���Ԧ��y�P����g�V�)ir�֏��9��W8 �+N�����p���U�y�$�~�c>��	���5V�����B�n=��O���$/�W�&Nꊓ�Hb�Tw���v�R��o�����F2]�J8�~�&T�S�F#���	���z�IYLy0�q��������H .�����F2]�J8�~�&T�S�:��b�>6"�F_hHbJ�02�@(]"Ke�����ڳ�/��F�Z�*�Rw�|E��L������8"_��o�߭�&HH�u��>��t��Vqx	��V�S����-ӻ�'4M���/=�B��YX�>� =&d=��O��b2�M/��J{K����Թ�4��=4���Tv��t�c�����Ä��V.�˸��"r*B
�	�`V�f�Bɽ�*<efMT�Ҁ����T�O����#���
�_d�Ǹ��;��2��:7P�7ٝGy��v��,��j`▘9���~
�l��������-�>G~ ���nj;T�v��S���*R	��Qo�X��<_"ƹ;h <�t-*��k�(�����ȉ=���$<+[�v������
���'�7� �EH�S����{"|:��lw�F_hHbJ��LD�r?���F1͝k���,(n����a1��F�}6�"��X��E$Jȝt�lL��Q�}��k���$��;j7�R�7��vu:׈S�y|��5�L/%r��^2D�"|�����E_�ֵb+�@�JПE�[5(`<��"$���1������8"_��o��hn��~���nj;T�v��S���l �R�|�����E_��VC}�R�)�+j�9:GA�y�y�����f�{��t��
�9����'4M���/�V�W�v#@5L�;�HrC{ѕ5��l��rɰ���k���,(n���M�����ӆ�澮/�žC��ky�-�뷱�nj;T�v��S����$4�ZsA�Y��g��<��ݭ�<����9�6��xx���]L�E�i{ޝ��i�t��Vqx	��V�S��F��q��v69k��8�↮GX\��М}��(H��u�6���ƌW�9�A���/^$�<U�������2�[ɽ�*<e؁̅5*'y^P%-H���}���)|�����E_��_��˴^�*^�XG>N�����·i{ޝ��i�t��Vqx	��V�S��@��������X�:��Թ�4��=4���T��, I!w�ɽ�*<e�+�r��y�f�{��t��
�9����C��ଡ଼�F2]�J8������MPⅣ�� ��	���A$�H�q)���	��[�bi�ܛ�|�$�䠢O)X:�?�^	%�
��nEbU�����|����с�*��2Z(��{:�?�^	%ͤ����lu�4�*+ZX��^�P��}��Pj�:�.��D��~���Cw�π[0H�q�DL/�,( 9������mr��%~���#�� (V���K��S�h��]L�0���{�(h;������7�dEe��?������8"_��o�������WLg#�^�F��������}RiY�;
��l�g!k]�:�����X��E$J��N��z�$��"�w��-�����yL�����"*����n4C)�&꺉Y4�:�M�Z���x�]�]�X$m2���jJRc�/u3~�l�QB�-�831� C��%�y<QP��򓤣�P1޸�.G���r�&�M��)�_h�l��q������f
� ���_ھi��͗
�rcq� ng�:�M�Z��K��
BL�^5)���ŕI�(^�;�S�ҚY
�[*:��:���N�	�.P�Ur���2�g�f�j� k����>щl����OX���(�D! �9��^��d?�E��- �.�Qq�*����p��݆=��'];��[0���߰�B��*��2Zڸ_��OifMT�Ҁ���%���K�z�6|"��K�Uxxb��m��Fo�l�ړ��ܧ���rzM=��`V�f�B'+G	�\ο�$Q����x���]L�EMͿ���q�
��nEE�(d��{E�6��h#A�Y��g��<��ݭ�`V�f�Bɽ�*<ec®p"�.��Pˢ�
x|Q��z_xZ��C�'+G	�\ΖF_hHbJ�
f�8�� "�����Ո�Ú�ȩ�F�(Uo��f�,+��:��:����mK�գ�������,4���?wd�ru��|�����E_v,�[sG��R�6W�m�R�5������*�-�_�av"�U��]��&����V2��	�G��a3I,�'W��VG�g~#��<�n�\��h��Nɽ�*<e�K�Sqr'
�R��ۓyP��OC��IǄ�s�ȠsoEu9U�s����Op�ű�Oo � Ѕ�g��e�ˎ�O��'���[���*�o�4ԽJ8<l������|�0E��Zɽ�*<e����M���4��]Q��x���]L�Eɽ�*<e�	������[�[]�ƣ_۫c����-�8wɽ�*<e�Y�tѥE�4�g T?0���{�(�rI��u��ޛfe�^C�ɽ�*<ekwO�&뿃��0ך��?r��U�e��H
E#LPA�Y��gu:׈S�y|��5�L/%f�{��t���8t��0.d�չ�R�l�VUQ�F2]�J8�F2]�J8�HE��޻',��~�� ��z_C=��H%zw�l�VUQ�F2]�J8�F2]�J8����D�dz�prpγd&[�ߌ�A���Uxz������Ą�#��MͿ���q��/�]� �V<\[82}5���P=�?�K��)�<�;:2��ؙH���/�]� !�d�`�I�v��,��j`▘9�ڭ�ܥ����k��-�)>˜y/;�)%��b0�~4�ɔ�ݲ������f
� ���_ޛfe�^C�ɽ�*<eE���7=��C�Ȩ_������w3_xZ��C�r�֏��9��W8 �+N�����p���{�m�f ����g��-V���z�]�H����jHi��}����6*HJY%q>{И��Cni�'\�g���KP0�>ɽ�*<e�#b����>&[�ߌ�(�k�$�0H��r�dZ�ŕI�(^��^����jHi��O�4��\"ɽ�*<e�YwVϛ��Q����_�'1QC\����2cm�Ӗc��<��^�QW�� �.�Qq�*����p����8t����/�]� ��ī|���^5)��u:׈S�y�է '���C}�/��cF2]�J8�F2]�J8�&���y���I�/K�P�;Z�F�Aܘ��'v�o.T\ۚ���h�C��ଡ଼�F2]�J8�F2]�J8��v�������2cm��d�p�6 }m!�d�`�I�NH���9�X��S�q��X�B
��ֈ2t����`V�f�B{��<Ia���� 3��;x�J�u�CKxP�:���X$m2�����UO`T�9���9��e�g�Q����_&y�AW>	ב���#m��)/�zC�~����0@��n�h� 	�%���K�z�6|"��K|�d&C�M��)�atBҷ��c A�[f��ԣ*P�k���,(n�|�2<sq�l�Z)^��_�������YwVϛ��<u��rnN�-���N:�r��NSad����r���)/�zC�~M�3pI^C��&Nꊓ�HL�"۠��JПE�[5'$��R��e�ũb�\�GeE+�O��N��S%��?T ]d��fo��ޔ�e�8����6+����E�	ah����ó�Ł#S�svs��
�������;ǚ J��B�����,(Q'ƽ���� �"�_엘������_�ھi��͗
�&�|�D��D/���z�<+��A�Y��gwp���	fH�b���AVDL��Lɽ�*<e��H7
kH��N��S%���
:��{gP�7ٝGy��v��,��}Rk!��^�(
P����|�1�ʢ:Y�f�H3UU���f�O@g�IFS�w�s@�����4�
�����%nġCB�I�t�`H�Q����U�xl�(T�W#�(�*� �.6p@�*3d�#_�0!s�,�	���
6�.8�0�T��(�H���-)�|�d!d�H�d�h�ݔ�x��{��õv�̟��������.s����g ��$�L��ow(7ALۗ)��/��	`�)�h��{̠����Lʉ/[¶���`���c��� �	[�w:���ע��������t��E�̎����D�<L}ڈ�����dn'y&���3��ͨL���K��a9q;���]��e�G<���ߤ#����ө�((|�w��M{� C<�ls���|����䋇�æ��tg������a��4W}����Y[A`�_Z_MyV<tn�||oKװE��"
8��o���l��͡U�R�4�t���#,�>�Y����,�:�+[��epՈI��	n��WO�.�<8��]���f8��H�\J����K=҉7�#������g~�nR�&x��l���Hwa_i��\{��ЍM�Cʌ���H�v���5������A��\��G������Oc]����s��� �F��.�8X��)8�\/,AܥЍ�ө�	I�\���YVeX���V�E{�49��������4�=z��F		DAu��6YhzoC-x�i���
V�r&A�V�6�.j���|R��Ǥ_�|�P��L���Xj��)�*��e/6�5��0�K(8 �%D\������A���UJ�l�t�p,|4�^,e�I��ހVh��)��&�I��J�ѹw���[�<,]�ͻlU����\�IFⳮ3f�d%\1ͤ9�mD�*cA��2p[�������Ɯ�h�Z��g)/x�*B��0�ѡlv���tk���I���v�D�t*�gc�꺉�@jB��Z�!�W�/�Cd�سy�%�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�]^�h��NI���}�N^���^��ˤm|���1f
�om��|G0�6��`ԬΈ��8��.��{�0F�d=R��蠍Q3MƇ%�u�邂�m\Y&�<��Zi?6�{�b��2[t�/7�`�$����-N��|��p�yJ���#a��}��V��h�Y�E��Rۇ�d=�����|�L��5:;�3-�Q��ݱl��j��!��}w���m��Z:S��]��\>�ﺚA�����j���7}_p��C����S�D��Ō�	�׿m~�,��o�A&Cr�,ԣ�؟�Z�Y�]��K-"�tI{����0����
����؟�Z�Y�'V ��Y��1$�g�P�q��{ȋ	,W�G���{�q�i2��л\7r����pK�ӷw����+���6���0����
���9s^���P�����%����%��!w�%�%ݹ����B�{��V�ڦ�<}"�22]���e�}��Y�Ru�"/}NzQBd���?���s�D{���]�6��b�X�G잠y��vgnկ�cm�/�8��w��e��(�iK�J/x��8��ჳIy�PB@����
�K����Yd�d�pqAdD��Ō�	7#�6�`��΁� M�#�|w+�n��i�  �=񣖗�3���{�tr/թ��A%o���:�\#����r���� fw�=��od��p�b����}����"��*V���1�+2��T�M-�Y ݧW��jh�D�F������dN���WI�r;�r�Z�����/|�T���fb%�î���}#��ha�0*�`�1~��7��q���TI�*�}\��C�>��������6��?g�w�j�hH=funq����>,��t���cU��w������j]�8�)I�&<@
�;ޖ�h]�7�b���DH%L��Z�âNxL �?f���8����1n���(!�8
�CB¬)<����0�By6JI�|�&;�
X�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8����T%�g')l`�A�I��z�gg+@1�H��;N
RC h�4�ZC%�45ԛ��}�6q75r�=�5�}�'ҺZ�ØK�^j����}��$EB<bb��i��<�a�]��S����a=?���X�t�K3h.���#��V�>Ey�U#�ɽ�*<e�M+DW��Ԯ�I��.��$(�dL	��D2��*�������%�B��=��@� �ɽ�*<e��~^-C���cW�e�>��9�B��K�ɽ�*<e"-w��-t�K3h.������L�� �G?�L��ɽ�*<e{*o��^Ԯ�I��.�Δ��B���fVA�0 y��*�������%b(X(i��5E^�X,6�ɽ�*<e��~^-C���cW�-�]�x�r8��6ɽ�*<e"-w��-t�K3h.��{`is3Z� �G?�L��ɽ�*<e{*o��^Ԯ�I��.�#"܇a��'~]�����*�������%Cü���8#.�E>2�<Uɽ�*<e��~^-C���cW��h���*b���]iLɽ�*<eEhJ9�һ�Fb�T�hAU6]?���,	4ɽ�*<e�N{}��ʘk�Ȉ�w�fx/#��0((�;̃{����a�s�f�"��� A�(�J!����;ɽ�*<eɽ�*<eHw^���*�}�{�'�]dv��ɽ�*<er���4GH�U�S$JsC��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�M��X�{��ms��u�,*����8E,��l-����*�}Pb~J�Hþ+��EB�)d����n��r�B���_5��3��F��;���,4���?wX�1�{��F2]�J8�F2]�J8�F2]�J8�$�䠢O)X7�+a$@)�v�Jɽ�*<eɽ�*<e�d8E��,-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q�ݗ	�[!_��H/z��Y�8��X�ƆE{��H �����A��Y�ư$�}����������n��r\#����r���c-֙k�����d˫r���_;8Wtw~�b���V���()�^�5��K+9a7�Wx;?xԖ߷w-CHv@�����)!)gP\�x*ّ�9 ���.�{���*B����@HW�x+t�W ��+�eN�@�� ,2!��Yr5Kd߂�
F{<��)�w��o쳰�y�6Y���Һ������t�A�����s��R��;�6.d1��Q�wN���&a��y��˾�Iy��*�ӭ��0Hv@�����)!)gP\�s�K��Y����D3���K�z굂��OI�k/?��ƪ���x�N����%.v��=<�K8#���j��p)��+�n�����'�K����}�0�i��Ƒ��$E�0F=ӻ��V����>Jz0���^ưVx}�)�R)@^��h�G�=��|76�A���z�%�׬�ĺ{��A ���r���G�ae����  I·`���|�B�	�
�s��Y",��K;G�����WߋW��zJ0�w,4���?w�ɬ���A���D3���K�z굂aNR̜v]�2�FF
���r����yg�ڥ��Hv@�����)!)gP\�.� �����x�z往��(���̈́����$ݫ�tF�ō�`�ێx�V����n��rF2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^f���!XkU�*�ǡ����QPP(,��*��:�mc*�D��|F2]�J8�F2]�J8�F2]�J8�F2]�J8�T�N�:Y�?���K�5߮ݵZ�?�	��$��h�>��@sy����+��	�l�M��1@~���$��| 5v�R��r��W��=S��jt[�n�>�Z��X�&��p��	��o������F2]�J8�F2]�J8�F2]�J8�F2]�J8��l��q��;DN-kh���u���@Eݟ-�n���*[���h�tMӘFʍ���{�_�)����Vo���JPAb���x#����n��rF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��l��q���{��ê�A�e7@(��a���0�&7Y�0Y�\��b��%L��V�81,4���?w1Z�w��1Ƌd#�a�VT���$���Ǵ9�A ��M���߂���T������a7�k��<��nG*�lۘ�>����O&�C�;:_���L�}�A᝞�����n��rF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��l��q�"�o(�E�:ɽ�*<eɽ�*<e�����&�\u�bn�z�X�1�{��F2]�J8�����q��XF�P��V���/��l�VUQ�F2]�J8�F2]�J8����IE/UeB^��r�a->�d��`�Âx>C}�/��cF2]�J8�F2]�J8�&���y�����:_����-���vGF2]�J8�F2]�J8�U����@�5����_k`ɽ�*<eɽ�*<eɽ�*<e�S����� ���	/�yl2����m�}�4e�YJ�D`�����)-:E��0{�I�n �u�HY�K��^��e��|>R}9��T�F-�U3^:j���+�J�DX�>H'����a->�d�wo�	h�[ɽ�*<eɽ�*<e�%,!u�r�"U�8?1A��!�(I�=LU[$"\�I;���ɽ�*<eɽ�*<eɽ�*<e3�lp���|M��t+cs��7Z���W<:Kɽ�*<eɽ�*<eɽ�*<ep�L�u*���I>/�4	�߅|��d72L%hQQ�J�1[�q��� E��w}���H�.}�0/+��=��c��v���W<:K_�������_M���5��^7�����Si���K�=�Zr%������l�*�[��^Us&v�%+XfZ�|�C��i�.�!/A�h���f����N���6����=�ɽ�*<eɽ�*<e2vr��{�j�s|Oݽ㓤F����Zr%��������a3mɽ�*<eɽ�*<e�%,!u�r���*�jCe�V8��+ ZH�ڸ��P��B�a�h�ɽ�*<eɽ�*<e �jv�5�=�̌L�+$r{@ �P�G�����F2]�J8�~�&T�S�F#���	�>)[�4�KeC��ଡ଼�F2]�J8�F2]�J8��a->�d�wo�	h�[ɽ�*<eɽ�*<e�P�O�_�	�y{I�7���k�L����z A�aiUj)��}w�u��V|ɽ�*<e�$��U�_���#��g�^�yl2�����h�����V��H�f����:��$��iaK�sB9Hl�+s�A�h���f��� ��#*ɽ�*<eɽ�*<eɽ�*<e�,8�(\��؊��SV8��+ ZH�ڸ��P��B�a�h�ɽ�*<eɽ�*<eȩ�Ļ�����d,����<���^���f�U��72L%hQQ��p��u��dɽ�*<eɽ�*<el<��b��x����Q���Zr%��������a3mɽ�*<eɽ�*<e�P�O�_d��ٰ#s`��S��72L%hQQ��	T(ܲ��~>�� j��Y��`�)��e�LU�yN�F�8I����N���Ϯ���O�>R}9��T�F-�U3^�G�3̣��[���MĞ�l�A�B�Z�����9��ɽ�*<eɽ�*<evS+ё@|���˨mG5�td'P�TT�I����N���6����=�ɽ�*<eɽ�*<e�G�3̣�����v��{s��7Z��~��Wɽ�*<eɽ�*<eɽ�*<e�]�F]������.�NH�Sk�𷉋5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8��AP~�;��jL���$gn�й���*�D��|F2]�J8�F2]�J8�F2]�J8�F2]�J8����.��Zݪ+i�uq��Xx0
����.o`�� �P1sGL�)��%`�� �P1sb����/�k��S�1�g:�.�U�[�Fux��z�,U�n[��p�rD�_f>�W����Qц���L��۬����:݌Zݪ+i�?�7��5�i��#SQ��K[�k���������t
Hp��u"-5�m�K�Zݪ+iG+��q�a:��`�8��:9y����HQ���y{`is3Z˨��ҮE=c@�LT'@(f]���
'��Ix����1-/gBem�]_Bs����LPnr����ˣ�+�����Δ��B���g�Xy�6%���Nbq�wԤ�ٔ����:94�+MO���tPfW�������F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�&���y�������&���͝�b�\3����ѽi�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�k��S�1����Ay�߿9�P��4wϷ�'�/E��Δ��B����PV~?�ow����@��Lsș����e�A�X����T���D�Cy�߿9�`]�#�ͥZ�4�?�C}�/��c(�|���
4�^�6�r{T-�(�|��3��]�����|��j�G����.X9ش1O�r�rz��4!���B_�h���*bk��xZw�~�L����Kbv�U+}�JYw�8�r�rz��^��tpx�B���tD�_f>�W����Q�/��~���@�X��?k; ��<:��u�;җ����V�C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�HE��޻'����̲�1{�:;�����R0;��L+�&�<�C��x�F��Mb��aO��q�I����e��Ƚ�L��F�W�����F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����%���&ꬶ�Rɽ�*<e�يHc~��F��T�l���!Z�_�'�=�3��&ꬶ�Rɽ�*<e�يHc~��Y���p�P��O���.��I@T��H!��R���e�DN
4��Y���b�6��۰�74�����RKD�vQFɽ�*<eɽ�*<e.f@į~����)O#�o����÷�L���
>i�]́�>T����>!�}����U��6���yߒ��`�g@�ȃwg��SY�h�/��I�04wݺ+5�*N�s�$(�dT�F-�U3^G�Y)S+�-}��5~��v����ɽ�*<eɽ�*<e	t�+������nX����ar��Z�.ɽ�*<eɽ�*<eWZIN���q._�+�8�zN�����ɽ�*<e�p\�Ì�G���.����сɽ�*<eɽ�*<eVG�X�y�k��٨S2�k-1�>l��Z������ɽ�*<e���Af/_.�*�f��vU�����_b�\j��ar��Z�.ɽ�*<eɽ�*<e��3�y���v�7��s�Z�����J��=x���zN�����ɽ�*<e�p\�Ì�c�9U�HK�ӈQQ��D�Y��3��g� �	�pm���Z������ɽ�*<e���Af/_.�*�fĳ�Ub9��Q�ͣZv�8�0ف����^�P��k2�G�Cz+P3�/���++����zA����%`�.�CD.�@�2�(��!�kΗ��U�I|�G�1�!�fiW�'"u��j�8]������g�g1�!�fi8>Rn���0H��r�dZ��<��ݭd��PtD��n�H��46��,\�܅�PZ���#dJ)f;��W��*3ZC�q�����w��l^��4^�Wd���U���������F���
��
�������%n��'����0.d�չ�R�;��f#Y���L*�D��|F2]�J8�F2]�J8�F2]�J8�F2]�J8�HE��޻',��.�@Q�Z�V��Kn��5Lͱ!���n�I���W)�"��|� -uR��Eo����b]qGt�s�p�LQH���P��%�AО��j)X�LOzyָ�˫�9�ʲ�7��&�UK} �l���Ģ�����&���g�w�6�+5�K��%2���L�-C�������k&��c����tn�~���FS��א�-Kc�3���lm��)��Rf�&���[ktR�/��Fs'�X�1�{��F2]�J8�F2]�J8�F2]�J8�	C7��3�^Xƻ�2��gƧ)�������~�Ǿ�������zxrF�hc7_��y�<rO�I{�3�Jc�8�akwO�&뿃��ѻB�p��Yqi��C�x�\��	�y{I�7�T�1�G�J'�k�[�I�s|ִ!��İ��U���N;�E�&Nꊓ�HL�"۠����GB����)��AŎ�HP�*�8⑇٨S2�k����p��}��Pj������lאHh�q6 �S����Ǿ,GLY/'��ơ��'���ʎ/���-�k��,��Ǒ�V�3U� ��,�kd�/�@.f@į~����)O#�o��`�7.\�+�r��y�Q���'�}�ٔ^qt�����q�E����mV����� A�[f�矑��ӆ�澮/�žC���U�8�sl�Z)^��_������G�Y)S+���(�
1�9'�ژ`Nɽ�*<e�i�J2�k�J�J=����E��-"7�!ne*5��uf}�*]��x��F!���8�!�|����,�4 �.�Qq�*�w/��e�	x�a=���j;�����p��B�N���㮄�I7ة��Gl,B!-.ȧ-4=�k~j�Kh�}����U�r�s�ec`<�S������K�`A�Y��g�����r��f�af�w�U{�$n�����nX�����8t��0.d�չ�R*����n4C�}c�\���x�\�C'�K��w���]����9����*�g�Me ��:�*����n4CO�nu��MK���7�2P?{,��t�ؠ0v3>#"܇a��,(<S�`d�����Q��0YJ=���ʓ�O�>�P h�ayAj	�����V��#�سLn%�au�*����n4C��e�^��y���z��+d)w�ٳ_�a�d��L�8l�=K�r$�_�kt�5���� ����6��۰��6VN�9���B	�D�J�DX�>HB�\��L���%,!u�r����������`.}�%,!u�r�"U�8?1A��!�(I�=LU[$"p�L�u*��������^��F�����_��ӧ�v�ਚ�Dxţ�v*_g��ن�_�����P���vz}ͫ#f���A�Y��g�l�VUQ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q��7C�Xؕg�Lδ�k���TB$��,�=�����9���5��#^�{2#�*�D��|F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~E�L�J�zN�����ɽ�*<e�p\�Ì����FKr��<�WV
v��6����=�ɽ�*<eɽ�*<e�N�课G�\DԷ��J�2���C�sNq�0a�w�u��V|�W�Xr:Z$�_x�'���0͵�Fb���g�H��Ę�c��<ڇ{� ߂���m{��v].�A����p���j����_yqWXĲԷ��{����"��Ip�ёg�L.M�"��G�"@cy��8B`}��:%�q/$x䴼��Tɽ�*<e<��:�Q����_��=^rgw�ƝCG��σ 6Uɽ�*<e+4<�a.�W��u3��k����p��8��d}���DhY��F�-I�����ɽ�*<e�r_�g-�������Mh�;�q�9����p��_�@2z��\�kܥ��qU���������������V�uCM+�n�/�G�M`.ᕀPI߬H��}!�Lڜ3D>�d�ɽ�*<e���1�f7��Pm�ս�6��۰�ǊVgrwɽ�*<e?\��ܰ��eD��q�d ��#�݁W/���ɽ�*<e?\��ܰ����ʕ�N�课G3r��?��ɽ�*<e?\��ܰ�?��N.̹�
�B7 �x�/s� �ɽ�*<eJ횈�r�֏��9��W8 �+N�Z��rÝq��?ʌ�7KS��ɽ�*<eGi
��Cj���FKr��(��ժ�S�����>�����ɽ�*<e�����Q��
�B7 ��9�����7�Z���_x�'������p��}��Pj3�lp��ܩѥ����!)C�Q�&�T�2+��@u:׈S�y�է '������g�HC}�/��cF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^YG~fza_# �RR}1�l�VUQ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q��*d�IS��_M���5g��*Kv�dx�$fs���ö�#5*d�IS����)D����W/�p.�qjX�f����F+�m9K�A)�^U�ɽ�*<eɽ�*<e��(`u)]��_@��%���"������сɽ�*<eɽ�*<e�A��Ǽ�\�����O�^p=��A)�^U�ɽ�*<eɽ�*<e��(`u)]�I�i}����9�G��ɽ�*<ec�0�I7�ar��Z�.ɽ�*<eɽ�*<e�`�2W�d�P���vz}���9�G��ɽ�*<ec�0�I7���jJԔɽ�*<eɽ�*<em�/�lvq�-�DzA��q�f�v��������g
,�C˾�`,!�^�)�OTC�M>���e`���T��|�r[ĢTYܻ�Mλ�h���H�`��ʄ0��Ҡ.�!4�HM>���e`���T������ovL�zN�����ɽ�*<e�\�e�=l1�!�fil���RKD�vQFɽ�*<eɽ�*<eOzyָ�˫�S�L�v�{�'�c� ����сɽ�*<eɽ�*<e́�g�N��,h�y�&:���(�E��ar��Z�.ɽ�*<eɽ�*<e�[18˞*K��|I*�j3��a'�=�3��&ꬶ�Rɽ�*<e��_��l�Kk��4;���OC�I0s9�>��b�zN�����ɽ�*<e:j���+���"�5�(�$���k�Z������ɽ�*<e��#2M)�}�
���*���m��ɽ�*<eɽ�*<e� 7maH���;�/��<�WV
v�����b��� � �oCU@T��w�9��ִ�[��L�)�d��&?ΦW�Xr:Z$B�\��L���يHc~��h�C��A���l�,H_��(`u)]��_@��%��F�����_��ӧ�v�e�/�K�am@�^������W�Xr:Z$���`�u�S��_9I�A��Ǽ�K�	�҉�!Z�_�}��BD�����)<���/�B2�:J�Xƻ�2��?�]�U J����D3���kf3����mK�գ֓o�D�a}��	E��{q���,�͗�O��ĺ����Q�>���`܋���-ֽ��
:��{g�q�И�mJ��E|�m;(��Î�HX	4o�1v��1�����4��`紙�����Tוۏ�@�8�!��=-�Nn�F�{#�M�է '������g�He;_��f>�/�K�R����)O#�o�����r�������M�1����L���	c͛t�����̃6!x�����i��ͻH�m?�GU0.n��_���v��{9���h�J�l�VUQ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q��&�!���H9iO��~�L6��ˬ�r����L7bZX���M�9Z�v��od�;��4[@D�cG�C�|	�ΰWs��Mr���V�:����݄�����dN��^Lb����3=HǎX��9ަbq<.L^O����w�t�C���"E]�7��|
f��X۹J���A�EA�)Om3f��1�A{�ż����Ǟq<Q��b�m�3��2U�L�#�B�)W�;H#�p�!������V+��@I�h��A2�m:x� �M#ċ�{�(�Q�
3�������NQ6B�X5A�}��?��4���ĩ���x��x�FI�ii�<K?�f�8(�)o*�KK���_%S� �{�FRA������F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�ác��Y������Q�\#����r�����]�lB#�<	ݽ�$��U�_���~`��rXuu���I>/�4	��oY��J7�����K�am@��F鈌E��i�����^�3�AD��%�}��WԱ{�R��:IT���s��'�MV	��ex��6	���ĩ���`��5���ṥ �u��2;E������с;=��/��n�+�b�?>|
ϒ���'�=�3���G��B�%�:�wD�+�(�T	�k2�G�CzՌy�6��h��%�~�������x���]L�E(��Î�HX�X&�㶮Ze�7��-�$@�՛�O���zc��Ze�7��-�>�����u:׈S�y��L��Ԝ�x���]L�E(��Î�HX�X&�㶮Ze�7��-�$@�՛�Q�%�g"'�&Nꊓ�Hb�Tw��5�o��l �Rym�To� T�uїKk��4;���OC�I��2�,I�>Ze�7��-�$@�՛���t���.����T�38�!���䱊*�jCe�V8��+ Zq�Qy[�^Nt+�N�K�,h�y�&:P�<(Ϲ�󬡻 �����luf:S��]��m��'T�*2p5m��:S��]��vL8q����{�'�c� �0͵�Fb����q�EĄ�#�⑤ngF��)�N7ֵ����"!k~��bC�`�x��cM>���e`���T��\�0=����[?�1�!�fiQ�(�eP5A~��"#ɽ�*<e'�9O�V��]}�[V8�}�9��̱�>Գۖmlvq�-�D�,m���<qc�������0H��r�dZ3ƹq�nNsցt+�5%�j3��aھi��͗
��讛 ��Z�0[�3�\#����r���V~��WE�i;�������1��g�eGY��J�h��
�����+��� �,\�܅�P�j3��a��U���ߛ,h�y�&:~��"#ɽ�*<e'�9O�V��]}�[V8�}�9��̱�>Գۖmlvq�-�D�,m���<q,xX�u���Ɔ��"�����Q�3�T�y��q����lvq�-�D�,m���<q����� �'k\���3%�-�b�f}�
����!�7C	�M>���e`���T��:��c]u�!�,m^$cIF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�HE��޻'�߁��`t��ߌ�VIרx��y�|1�#�T��8>r?0����v{�1�N�-�(�[΂����\$�� f��5���i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q���~�>�p^�����%kw6�6�&�'4M���//�%
q�s��Kv�V��P1޸���$Q����x���]L�E3ƹq�nNs�]�|tֿk���,(nĐ��]}�[V8�}�9��̢`5V���A�Y��gV�������d�a��|��p��E��o��ɽ�*<eB�B/"��S�Ÿ,w%�y�[Zo����8�!�|����,�4 �.�Qq�*�`V�f�Bɽ�*<e�Z�0[�3�\#����r��_؊��\���,(���W��d�a�ցt+�5%�A�fɽ�*<ex�N����!*�,;E��O��]�Q�>ٞ�ć��}Gδ�-3�T�y��|��R���m�EfܰP<0�����Yr5�ݭI�ҍ��r0�w�S�<�G���u&4'�`��P�[n�b'5yW�/k�ۥ?M>���e`���T�Ϡlr|*�.�+�L�t>�L�������p��h��;�p��/BƷ?�yN��d3M6�3��,q��J.
�XC1��q�g��������H׭P�h���������|�{��"�p���U��ɽ�*<eǩ�m*M�5V�K��9��U���ߛ,h�y�&:�e��0.��tuA��s�,\�܅�P�j3��aھi��͗
~���y� �+)���;C�p�
�a>���`܋
�Ҭ��jQ���l�Ѩ�Z�����������3=�t��ɽ�*<e��p^�S_���N~�E&�ݪ� >��ߖ�Ilvq�-�D�,m���<q����� �����M�bsGj�{sN��8H�Ϸ�?{��)�w׽�P�7ٝGy��v��,���A)�^U��5f���ٓ�l藌V��DLfF�b�qU�ۜq�yf�_��#�{#�A)�^U���IG�P�����HZ��O���.���i-��4���ˎϱY�8���ለ�M^�0��%�~�������.�냼L�} ��y���,ߺ�z���;�V�2E}L��3 ����28:�������p����{v���G45Z�)��,����nX �q�ƛ>�_=R<4�=Y�,�����+ Ң�E��_��#�{#ɽ�*<e�}���O'�i�C#�Me��"ɑkH�E�s4�vZ'��v���g���-m�q�*.�k�Q��
���<�WV
v���d���t�Q�L<��_��l`t�c&�r���[18˞� ��R�>G���#H��i{ޝ��i�.�
�$���5-Qo�����Bg���4�2p*ۻ�9�A�Y��g�A)�^U�����!�dg�Ycw[_���[+���(l-)QoxcW�x��xA�Y��g�.U�[�x�G���H���������0�"��S�Ƃ��� ��ʅ\���%eس^�d9ɟd$���fg�2����p���ar��Z�.ɽ�*<eɽ�*<e�����3t�_=R<4�=f��{�j����g ه��V���P!����p����{v���G45Z�)yLk IlK7�����3t�_=R<4�=Y�,�����+ Ң�E�ȇ��U�Ԝm�.M{=�#S�R�L������V`A�s��VJUT���i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)Xɽ�*<eY�؟�r�C��0�� ��ʅ\�)�Ŀ1.'΀r�3�"����p���{nvC͎,4���?w�}�2��;cu-�!�J�
��?M+�`A�۶�D@7D��6-�����$�L�!&ǋ�E��,4���?w��݇%�G���h��nr�6��[RJ=�bL�.��	��B�fn=�D��@��6އm��U#�VJUT����{�;���R��蠍Q3��rlT��DGAR�ݯ�b��x��t����
:S��]��Q{��%ߕ��cW�Y[v�_�n;1D<��*�m^w����P�(�w�}&�����Rq�y5�§]�o5o���w����p��NM{9q�����y���{�������y�TAA��;}������n��rVyB���ݗ���㪯hgM��hZ;����|:l/����p�g#*V��L],'�P��ݟ�+,4���?w���چҝ���0����YK�Nf:+�7ڸ�3g��[��Ll&)./�"YM3�
!8�f5�I����,4���?wmP�����I�<� w*qoƅ��tu*��3�/�����6�~�������p��C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����p����{v����$(�d��,����n������+�8j,~��¹���ɽ�*<e�2���
�׍}JpE�I����~kf6A��-}��5~�����p��}��Pj�$��U�_�*�W��(����Z@,\v�n �u�HY{��\�jb��{�?����[��RԀm��P^ɽ�*<e��Yr5X/��m�9uERd�($
��1����,w¨�]Mg�4���9V��Jm2��w_313�����K�a=ɽ�*<eg�D#$?��(l-)QooW��$�O*(���4�6I7��O�M�b|�5�px�����������"�@���Ր(l-)Qo��0nҰ_�����p����e-���A]_2�\��EVkB�#I��.Gh��d��6��!�=4Y�
�u#f�.`��6�J�1���Jj�����ɽ�*<ep+��cۢ^p��'�K�Y��vs���JK�H��2h���76�^���e�h�ɽ�*<eh��]L�T��NuO�/����s������^V7�@3�w�~���I�ȝ�%1�M�@ ��:�����p��C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�M��X�{����5>�V����5u1_���׹���۫�{}�-�T9��4��"'H�ɽ�*<e�����F2]�J8�F2]�J8�F2]�J8�F2]�J8��l��q��A)�^U�����g
,�\�M4�04���jp�~�>��|��T�Ȁ6�,�~!�A�Y��g�A)�^U�����g
,��W�X�u3����k$���|��T�Ȁ6�,�~!�U����f��{�j�A�Y��g�A)�^U�����g
,�\�M4�04���jp�~�>��|��T�Ȁ6�,�~!��lۯ0�X{�kc�aSg��|��1"7�!ne*5_G%�1��M�H�D����Y��`Uaz)��I$jj��n��^ax{k�.c��\/�`�!:�~���6i�ɽ�*<e����Zɽ�*<eɽ�*<eԯ~�5MJ�ަ��[> ��.%��IG�P-C-h��P@p�y��`�7.\��^/a�Ͼ�2��t��;�+����l���*(���4�6I7��O,+�
����,w¨�]M�7BJ����9U����f��{�j��Ȝ����*�W��(辙^6v����j�8]��Q��a�03�3�_�_3��B����ɽ�*<e��*��� ��ʅ\���%eس^�X�t�.�D���S�cW�S��57r�<�܌���xy�ɽ�*<eG�爻>���F��,g����X�ڲ�
��@>�Q�?;C���u�̌�Wx�R$��"�V,�wda��(��؀�ffs�mU�p���a�o���Qtf�J��	��(ɽ�*<e���c٘p�ڇ
�܎[;��x;C��{�ϣX�v} �����a��fL��T���;ȊUܗɽ�*<e�;���n��`i2-� ���2����	��s��|�T��C�	���[Ϛ*ݭ�ƪy�Wi�u�R7�b]uQ�u�b|N[�
�	�vp8�$1���~.ی$�A)U>6�a?*�F޴#_��� ����A���a��L�0�)�w׽�O@����D �EJ(�X8Q����s��i�C#�Me��~�(�|��v�[\�ɽ�*<e7� �{�|�-�w�ѕ�"٦���7
���lm��*ǻ�F�kɽ�*<ekwO�&뿃�x$,��|��T��E�fx>�"Cg���b�B��EVkB�# �X���}1f�3S��	űQ�曔�g�`C��̹�`�7.\�ɽ�*<e}��Pj:S��]��ˏp�S���{T?(.�����$*�W��(� �X����龤BT��4����Ό�g�`C��̹�`�7.\�'$��R��e��Ȯo�z�ɽ�*<e�5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S�ɽ�*<e�;�z�n��f���d��x��j�flX�QE.%��A���C����ԫ�����*�~~��9§��V�O ����[Y�3z
����N� )qP(u�	��ݚ�	��ľ����|��p�^ֱ̾��d��-5�h(�(�| �����t%}��˰�$���x� ��ʅ\�;�R�1�*�7OX�bhiaI4�S�x>�{ȋ	,W�ɽ�*<e���V<}�OhI�ԍ��I�X4�YN�m�6��9��ڇ
�܎[�y�Sp����A������p��Vk�'r-׸��u|���Kb���*;\�]p�e���m��	�I��~G~�S_���M���|���!��s�biL�.`�))����)�Ŀ1.'k�R�F�y����8t��0��gq2q�R�sȝ�idRt-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�M��X�{���Q��L Ƶ8ׅ�$�}j�L�lI�Ml"TJ�\r���Y��q@�v-aDk���)���4b��&��F1����G$-?6��c�VJUT��ș�9����+�Nn��#��.�*��)��y�����G4u9<�������p����`,��T�VJUT��ȋN�h+�V�p*ۻ�9�	i+�����)*�Qyp*ۻ�9�r�,����vdi�xsIz�$�8`�;oj3[��M3)�$x�\�uɽ�*<eɽ�*<e/g�����qs�Pp�s�K��b��@e�'sȦ�Q%U��$$���̥H.����',4���?wɽ�*<eɽ�*<e��p^�S�"�h-P��|z���}O'��˼��1���0���Yr5�ď����1��|��T�Ȁ6�,�~!�������SZ��C�K0ɞ�BΉ�/@1��ϭ�L��|���E6��b;�S��BEtg]����"b�ɽ�*<e�����ɽ�*<e9<�b17�����	"�x�b�2�:%͏��ns�ů�C�K}`�Vj��Y���o���	��o�kK�ȹC���`�����|��T�Ȧ#k����*U��m<p*ۻ�9��uY'���-����� ?�}�س��v])�rtnFM����A)U>6�a?Y[v�_�ɽ�*<eɽ�*<eC��>�*\&kخ����%i�z��().11��w4���Za�G���Z�Jf��8��,�z��ɳ_t����>Nk����n��rɽ�*<eɽ�*<etE�6&��().11��ww���J.fG�%����(l-)Qoii�h��&F!g�x�\�uɽ�*<eɽ�*<eW�w*�7=� ��ʅ\���%eس^��,~��6���I��F��e����+�Z#hQ�;�+��gƧ)����Y[v�_�ɽ�*<eɽ�*<eu����fK��4\�g~1-o)"SIֲ�(���A�ڇ
�܎[��_�i�4�(��ј�>��Ȟ 2o�����n��rɽ�*<eɽ�*<eSNA���(�1��Ӫ*c��-C'2���/�9�1�ˮ��,��,w¨�]M����3�^>���e_U�VJUT���i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)Xɽ�*<e-|�V�P����A[���i�C#�Me��~�(�|�w��ﯢ��b<k��5MJ�ަ���+��R�*�&�X�Xɽ�*<e�T�t�g��g�����6��n��_Lq f�&�a�\C�Wd�ɽ�*<e�f��<j9D�m��ɽ�*<ex몋����U���Ɔ[E9錎�{�1��S�ɽ�*<e+�n�/�GcnNMG���뿓��'c%���n� � �5��<�Y��{66����)U�AI��"�׍Le�.�~f���[(�0F�d=������ɽ�*<e�}^B�Ņ5�{AM�ɽ�*<e�ޒ�Q�l�{����/�ӸP�[$z�MnhɆ�ɽ�*<e+�n�/�G>R}9�ܽA2�*PD7�3]N|�ɽ�*<eɽ�*<eM�Ń�����	/��-��)ӕy���V�uCMɽ�*<e4�e/.����B���R��bT�>A-��B��nɽ�*<eɽ�*<eo�d�BjZ@L�cs��U��h������p��ɽ�*<e�I_�I�O�Ph��Bf���d�M�.x^�p���ɽ�*<e<>�u�yo_��-ϓG*u����G�v=ɽ�*<eɽ�*<e��R�Mq��j�;�y	�^B�������cW�ɽ�*<e)� ֪w 1�@ͫ�����e�ʝ����ɽ�*<e+�n�/�G����Ph=��t��oGs���9=ɽ�*<eɽ�*<e�����΅���8�3���Yr5ɽ�*<eiT�F=U�>ɽ�*<e8��d}���DhY��F�1? ��6�5���@Ԁɽ�*<e!�T9���."1Do��CS�����d��V�pɽ�*<e+�n�/�GAiq��%ɽ�*<ex|�햻�E��%eس^�d9ɟd$���48"�It���cW�ɽ�*<eR㠍�������-��ƎAXU߮5MJ�ަ�����L`h��)����ɽ�*<e_�@2z��\�kܥ��qa�磅"��qi�r,��bɽ�*<eɽ�*<e�<�����49�iv (������7ψ�az�L����V��j�&�������}��[3��W������ɽ�*<eɽ�*<e,؏����q]�iʳ1�͉ ��ϗ�#o�yK���%/�JD'l��IG�P����aVl�v�W�-ɽ�*<eɽ�*<e�=X�Soj&��1��]�Nv��p�� ��R�>G��o�p�#L����p��ɽ�*<e���4\MP�m��"�,w#sAyA/��6����[ɽ�*<eɽ�*<ej	�%w\�����(Px�&Wɽ�*<e1C\ߜ��C�b�MP�+ �0��MK�s�Zɽ�*<eɽ�*<e,4���?w��=�wY�8�w ��ɽ�*<e+�n�/�G6���N%�&ꬶ�R-&J�� ɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�fɽ�*<eɽ�*<e���L��5�'��,��i=�Z ���ɽ�*<eɽ�*<eɽ�*<e��M�R��Lc �ھi��͗
ɽ�*<e!��(9�i���!�)�i���~F��mZ �/eJR�k�/eJR�k�/eJR�k����l�<�o�����/�\ȼ�]$=��ɽ�*<e�O�����X��Wo�������g�����l�ɽ�*<eɽ�*<e�VJUT���	D��:�^|�x�k�O�ɽ�*<eɽ�*<en���k��d���^���Ǘ����X��ɽ�*<eɽ�*<eɽ�*<e��M�R��Lc �ھi��͗
ɽ�*<eo�-ᛸG5�td'�tT���'%萚 tɽ�*<eɽ�*<e����n��r�����/�\ȼ�]$=��ɽ�*<e =s���GJ��tL:W������of-&J�� ɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�fɽ�*<eɽ�*<e0<^��`3��!�(I����-P��ɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ
��,�fM�ɽ�*<eg3�GIJ�"vЅ\�J3�W�`>+�h
�K=4ɽ�*<eɽ�*<e,4���?w��=�wY�8�w ��ɽ�*<e+�n�/�G,[h�
�+ɽ�*<e-&J�� ɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�fɽ�*<eɽ�*<e��U
r	]�'ZC���^1�?q�-ɽ�*<eɽ�*<eɽ�*<eu;�Qݷ�2U���m����p��ɽ�*<e��f`>T��u�d}l��{��Q�h
�K=4ɽ�*<eɽ�*<e)�,3u�A��e6�ڡ
��,�fM�ɽ�*<eg3�GIJD��ݹ�V����pɽ�*<eɽ�*<eɽ�*<ej	�%w\�����(Px�&Wɽ�*<e_�@2z����K�`�+ �0��MK�s�Zɽ�*<eɽ�*<e,4���?w��=�wY�8�w ��ɽ�*<e+�n�/�G)�7h����X���b��x���ɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�fɽ�*<eɽ�*<eJ횈���8t����"�z7��yΝ;]��
�;�+��b�Bo���ko�%����Yr5*�D��|F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^�VJUT���[�ҐcS%iv��;�3-�Q�4�DFnV��ꜧ��o��g�Eb���(�nf���()�^Qc�k�"u-�!�J���T��a�,\�����e*�D��|F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)Xɽ�*<e����q�E���蟣��B�3/���P1޸��\ͯ�R�ɽ�*<ex��*��~�������ɽ�*<e���U�8�sl�Z)^��_������ɽ�*<e����:#�3�3�_�_�qpe9|ʐ���L���ɽ�*<e�Y�tѥE��䅓�g ������ɽ�*<e��}Gδ�->���`܋
�Ҭ��jY�v�<�[����p��ɽ�*<e3����k$���|��T��$�ױ�ӵ� FsZ��b�;�+��)��J�B��?��W_�@v�zO��{���:By��{�&�(~�����I�z�(l-)Qo��9	�(+��
:��{gɽ�*<e��8t������p����8t�։0͵�Fb,4���?wX�1�{��F2]�J8�F2]�J8�F2]�J8�$�䠢O)Xɽ�*<eY�؟�r$�E<t���M�ٷ�O�6��SZs��cG�C�����p��C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�M��X�{���?�Vl��n]l� ����f���5<����]�DƄ��5MJ�ަ�B���)��u�i{ޝ��i�.�
�$���5-Qot��H;߾"
���lm����wEQ�K����p��]���/�޵[�Fux��E�I����P�o�|,`�A�GYK��,w¨�]M��5O�GLLɽ�*<e'o���.1��Be�5E�k&�r��ˮ��,��,w¨�]M��5O�GLLɽ�*<eh"J��aiUj)��}E�I�����S�Ƃ���;H#��J�~s��͌r�����?�Vl��n��h�������c���><�>֠�]��Zi()Ze�7��-��K�`A�Y��g�A)�^U�ɽ�*<eɽ�*<e�i{ޝ��iR�[Ɋ:�Z�ͥ�!���"������p���ar��Z�.ɽ�*<eɽ�*<e]��Zi()Ze�7��-�"vЅ\�-�f��ݬ"7�!ne*5�zN�����ɽ�*<eɽ�*<e;=��/��&�}��z&��\DԷ��J�VJUT���i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^�VJUT�����k5R��y�ƱJ4uG\$�uvo''w.e�������4�1�;A��B�,4���?w]^�,��7�U�H����u~�!�岫�] o���$��%����$B+K�,4���?wX�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q�ݷi{ޝ��iC?�zI�WE�I�����S�Ƃ���uQ���&�2��z�O�. ���vS+ё@�{.p�"��,����n���)-:E��;H#�&���r��8�d�	��ɽ�*<e(���|絪����*�ɽ�*<eJПE�[5ɽ�*<eo��^��;�I}Ǥn �u�HY ��A`��]C'�K��w�'�$j�ܑB9Hl�+s����U�e����T�LG5�td'd9�~����d,����<���^�0)�D�ɽ�*<e�+�r��y�����p��}��Pj�<�Q�E
���lm��)�Ŀ1.'Lf��PԢ��(l-)Qo��9	�(+5�3�4ˋ�K%J dl�{����/�ӸP�[$�7)p7O�z_*e"���|��T��I|��)5`0H��r�dZ(��Î�HXt6��y��]0p0P�t�(8.K�e|�;�+���;�����,+T0[��}5MJ�ަ�u�-^�Tv�(���Ww�fx/#��0((�;̃{���U��β�"ˮ��,��,w¨�]M�+QV�9�����-�8w�ל
ϙ� ���h3��M,�	���P1޸�l�Ik�yl�m��Fo�l��c��d6ɽ�*<eJПE�[5ɽ�*<eO�
�����GbY�%�JПE�[5ɽ�*<eɽ�*<e��f�仲�;�+���]l��+nL���L���ɽ�*<eʳw޿C�,+T0[��}5MJ�ަ�/�EL�Fe�NSad��ɽ�*<er�֏��9��W8 �+N�����p��ɽ�*<e3ƹq�nNso;t\�x���{|��SWq�Fd9@�����C����j;�����p��ɽ�*<e��
���(h![�o�2W.V}e����K�am@�Z`��'0頞Ks���A˃�6��Rb��fQ��;ɽ�*<eɽ�*<e<�D�z?����+�Z#hQ�;�+����F�n�]0p0P�t�(8.K�e|�;�+����޶(:ɽ�*<eɽ�*<eK������|��T�ȭ+2��KNP��]o���f�仲�;�+����޶(:ɽ�*<eɽ�*<e1��0ɽ�*<eu:׈S�y|��5�L/%ɽ�*<e�+�r��y�ɽ�*<e9Sz��l�MȁUN̩ׄ�$e��ɽ�*<e���4zm��QF��V��}�\#m^�~����p���c�xl{]��;���&wv��ȍ���u��-�/	�r��Q��FhvE$�y�Xk��Y|��:�'V~����x`��̫ɦZ�^y,4���?w	ȸ	^�6�����g��̬���l������+�~�`�/���M�)n!��~�0�7M#=sDJ7�{"]�y&��tt�
����h'ɽ�*<ex*ّ�9 �47*�8!flPӄSXWy�k4���nu�q:r�ط<26G΀��{2��V�Km��18l{'0+@[�VJ���E�ɽ�*<e���vE���`;���L�~���C�)���:��?�v�����D�����jܞ�̧��߉}O%� S������vğ�ɽ�*<e?T���׍���G�MR��o��|��ɽ�*<e�����Q�p*ۻ�9��[ŏݣ�C�p%m�:���IG�P-C-h��9ݝ����_=R<4�=Y�,�����+ Ң�E�ȇ��U�Ԝm�.M{=�#�[�fbKT��NuOrP�mW�(��Î�HX߯�d?'��v���p%m�:�+ Ң�E��fM���(ܔY���o��v���lr�f��{�j��lۯ0�X{�kc�aS����DǙK��WČ�  ����p��}��Pj� ��ʅ\���%eس^�"��`=����Jg�W��v���dLf�2N�2��,+�
����,w¨�]M�7BJ����9=�D�VtrT��NuOrP�mW�,4���?wO���U��2�Hq�c{�cb�}���p*ۻ�9�"Y���-�k�1I�<�ò�K�	� @�� 
����Op�űҍ�)�T�<Ɍ��;%P�����d��@Q=�n ����n��r����un!2�&�f����S/�����oZi#���q������@1g�eJ����Ѳ����(c���3�cdV��F$%��i�;���������kV���()�^׃"�|�(��w����9�k Y��w_313��8�)I�&,x<+d3�-C�������1و�d��E�[�ԏ�����wa�kdk�r�kwO�&뿃:�Uez�|��t�� }Y/�Q��N���!X�'��-Xpu��/Yw��6�#| �+*,+�
���Ç[3���pa�T	ʪs4z�3��gⴼXA5%
��=A&� ��ʅ\���%eس^�"��`=����Jg�W��v���dL�+�(�T	�ɽ�*<e����p��C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�M��X�{��N����<�B�=xyxNm�t*^x��ύ��>�����p��C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�M��X�{��P&�'s�G���0��(#�%X?�������~b��i���sX!�����p��䴼��Tɽ�*<ej��_h�-?�1�p%�F�����a���V�uCMɽ�*<e�-[z x�`���P1� ���\h88���cW�ɽ�*<em&Z��f�ӥB]��tFVd
P���kB��ɽ�*<e��x<�"l&�����w��&`!�D�_f>�W����Qї]���u��ɽ�*<ej��_h�-?�68�Fx��,D�qi�#-�g�sɽ�*<e�>�|�Y�R�[Ɋ:�\_:7�5ɽ�*<e�\	7Rn+ɽ�*<e+�n�/�G���Xv�k1? ��6�5���@Ԁɽ�*<e�r_�g-�������Mh�se�gې��h
�K=4ɽ�*<e����p��ɽ�*<e���1�f72��S@�`��uQ���&�2��z�DS&63��ɽ�*<e+�n�/�G�M`.ᕅ��~�I���깱c݁W/���ɽ�*<e+�n�/�G�F�W�����CS���R�[Ɋ:�R�S��� ���cW�ɽ�*<e���!������b��M&��hx_� &���r��1vdf�f�ɽ�*<eɽ�*<e?+�o&[����2c�I���ĩ���`��5��h
�K=4ɽ�*<e����p��ɽ�*<e���c�=,�ӻ��)��e�LUW:�=����ɽ�*<e�)�w׽�ɽ�*<e��vVK�`�|�` ��"�.�!K
5MJ�ަ�H�M.LD�~���cW�ɽ�*<e�Ll	d	�zRG];WJ�\i:5,w¨�]M뺽�7��ɽ�*<eG��.s�xɽ�*<e�j��?��8ɽ�*<e�����F2]�J8�F2]�J8�F2]�J8�F2]�J8��l��q���MB7\]P��X��[�~
J��A�ύ��>�����p��C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�M��X�{����^/a����{^X�G�Oa��Dmwj�e�R�[Ɋ:�}�a;4�����hBx�g�+��'��)D����t7v�H�����p��}��Pj�;H#�������cҘ�]Y[�P���ĩ����y�\���R��'rr~�L���:�%���{_E��a���_ɽ�*<e�
���ji����ĩ���F���YV8��+ Zjbu}�^�n�+�b�?6�3n<q�$V �0��j�8]��ߒY	T�%�:�wD˃�6��Rb.���\R�[Ɋ:�}�a;4��I뒒����ɽ�*<e�����F2]�J8�F2]�J8�F2]�J8�F2]�J8��l��q�N7h��IkGq,w�M5	�6���5E���E�Rģ�t+������n��r��&���6����v�M�[	�Q��ԡ���,E�E��2�~tAt�VJUT���i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�~�&T�S�ɽ�*<e��v��~��Q�YC��/�žC:j���+��&�P����b��M&��*���W�Xr:Z$O�. ���ɽ�*<e�G�3̣��l>j�m�ɽ�*<e=�PM���%�:�wD�+�(�T	�ɽ�*<e�]�F]��Ф����7ɽ�*<e��b���Ze�7��-8�d�	��ɽ�*<e�]�F]��н��g�@P�G�c�т��b���Ze�7��-��K�`A�Y��gȩ�Ļ���̢���k�!�(I��SFt�aWq�Fd9@��G�N2�Wm�B���p���b�!�vS+ё@_�`/I�W6���<���^�w�T��]��;H#�|����V8��+ ZA�Y��g,4���?wX�1�{��F2]�J8�F2]�J8�F2]�J8�$�䠢O)Xɽ�*<ePk�����x��q�k�gΐ�Me���=t�rt������ܷ���I�%���dN�=<�K8#��ɽ�*<eOpix�����Ds��37��ڜ�ɾXe�g:!�'R��ɽ�*<e�����F2]�J8�F2]�J8�F2]�J8�F2]�J8��l��q�ȩ�Ļ�ԁ�uz���d��-QJ��b���Ze�7��-b:n\����2Y	���FD#�����z��R�讎��yK#*bt��Oh�28�;��%�	X5�Ӿ��I/k �u+�%0ɽ�*<eU�����gU�*�ǡ��^�Ԙ4+ޛfe�^C�ɽ�*<e:j���+��&�P��t�ؠ0v3>#nZ~�n�4L}A�\!����ɽ�*<e�)�w׽�ɽ�*<eO�
������*g��-���Ծ��#��V��@��S�>�-�ǖ��(��ս�@�m�##����asE� �v�x�|fh�*�&�<$�9�n��Y�hE�	_�u�n�`V�f�Bɽ�*<eɽ�*<e�>�pؼ&��N����@z�Jɽ�*<eɽ�*<e�$��U�_��ѥ�����O�pٺe�ɽ�*<e'$��R��e�����kV�'$��R��e�����kV�T��%z�@�(�=ā~�"��}��u:׈S�y�:�Q��d[�k�s��٨S2�k�8ߜ�R��������;���
N�Q��s�B��{����/ַw��g�.S����YT�F2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^��ԅ?����m>�u-�!�J����}�u��볯`A�Ɗ����F2]�J8�F2]�J8�F2]�J8�F2]�J8� �y�V�����tQ<[f���D`��`V�f�Bɽ�*<e.}�0/+�,�o��vɽ�*<e!)C�Q�&��K�`A�Y��gp�L�u*���L�PlC�V8��+ Z. (���9�p_�>oXm�B���p���b�!��0{�I�+��%�ٰ���˫񷗤Vk"����N[�V8��+ ZA�Y��g�_פU�/�%�7㫙�H���8M�C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�HE��޻'�S��ō0�<�>��*�Eo%mFi��>��(�Y�,W�/�5�|��}\W1'4�X'ĳ��adg�Qt������F2]�J8�F2]�J8�F2]�J8�F2]�J8��6(�
r4�w��g�.S��}Gδ�-�	�=7�PsC3���c{�j9������#���),�߫��Dan`V�"�_�ɽ�*<e��v��~��Q�YC��/�žC:j���+��&�P����b��M&��*���W�Xr:Z$O�. ���ɽ�*<eiG��?\�9�,���Xe���g�Qt�ɽ�*<e�G�3̣��l>j�m�ɽ�*<e�,S1�;��}!�Lڜ1RMQ¥�ɽ�*<e�)��e�LU�!I�2ɽ�*<e�ew��7��s~;fT����p���P�O�_i�.�!/�B�"���p��u։��2��z�݁��!8����p���P�O�_!`h FH�
�̸B���a��b�*��2��z������d<���J�ܰ�rɽ�*<e�]�F]��С�W���#��U��Z����ܤ�J7�����K�am@�p���b�!��VJUT���i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�~�&T�S�ɽ�*<e�/�����P�
�XPYp���ل����|�L��5:��8���6����O�
f+��njiɽ�*<eWA�fV�����=(�/u�� u�o�NQ�sK��<k#Sɽ�*<eC��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�M��X�{��vS+ё@�2��z��5����)��e�LU�ܞca.o������/������� '_��~�Z����O��B��l�iV E��{Gɽ�*<eU�����gU�*�ǡ��^�Ԙ4+ޛfe�^C�ɽ�*<e:j���+��&�P��t�ؠ0v3>#nZ~�n�4L}AEu;��%r�ɽ�*<e��
�����?�@ە���F���
��
���
EÎe?��zk=��=:.�[�r!w�iϞ��Y�hEK��|А]zI�v;�8i	�
�s��Y",��K1�w�w1l�XiI�����p��ɽ�*<e�]�F]��о�~-y7�A��K������p��ɽ�*<e�]�F]����I>/�4	���7�quA�Y��gɽ�*<e�+�r��y�ɽ�*<e�+�r��y�u:׈S�y���|�r�	~���&Nꊓ�Hg���J@x h���2&/1���	D�ܣ{U/��A:��i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�HE��޻'Y ݧW��j��0����7��Ѱ�iXm=�4�i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�HE��޻'���q�����T+8!{,�=��aOFP�
��ߤ�y)�<zeO�sΉ��WxBW+K��⳦@�v-aDk�kخ���v�s�ɀ�b
������.ล���3�<\��S�8��5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�00��[n���X��X����
����Aę%���<�2k�G�d��PtD���lVܜ�������9PG�2���(��Î�HX�Iҗ��n�?�m�v�֜4�r̎��`[�"�o(�E�:�X��f��Sz�AO(1�!�fi�uTJ���i/�{lM>���e��0o#�����Yr5ɽ�*<eɽ�*<eɽ�*<e�S�<=����S�j孖�Y���m�V�%�����D3���kf3���˪�%�&���z���z�7T�S	L�v+��i�T��%zؕ��g�q\���%#骜NעD)������?5�j�8]��O�j�<��ֲi9��i&�:��@2�<�_xZ��C�����,�4����0b��*��-`������F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8����U����!A:����i�2���4ق�,���)��b�d �E����!§�v*"H+��b:!�'R����0�Ře<I�h��A2Ƙ�C��m"��O�+���D3������8j���A����N���d*���݄8�n���"�,���)��=�$lX);�3-�Q�TIIK��<��ҵ�C��?<'8D��s$|��C�p�GES(=lbP���]�����yU��.$����K��7��P5L�ЗU%?:��>��W��z�[(�gԸ�N����" �#���t�R}�n�c3��Γ���)��Hv*�D��|F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F���3��ބX��X����
�������:^�H2S鋅$z��Áu8��l)���O�ة�w��ɽ�*<e�����Q��5f���>}�e�Yw�\�%�%�L�'�����H�d��1����Zts�2� �������|�{��"�2>Ѭl-��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<ej�`	n�[�I�i}�xh?��60��JZv�W`J�#��P�� �>�/~-�7KDd�֦#�[��޷-�E��A�Y��g��<��ݭd��PtD��N��|�ISi���E�W����p��}��Pj�v�s�ɀ��O���.�ƺB�9�IC���m�ö�������᷻0
�QEo%m5��#z�^�c�9U�HF�Jf#Գ��F#���&D�� �4~��o���!��3��֪��	D�ܣ{U]	ȳ�ؾ�k2�G�CzӇG����!rre�N�� NO�Y@�ܧ�WG�ӌn�U�{�"	y�r/u����v���b��
8uVT?a5Kcɽ�*<e�����Q��5f���>}�e�Yw*��>���>�D�'�8���`��FG$;^5�� �	���{���u�P�Q٥���"��m¾�H�Q3����Lc�k{�sE� �v̗v�s�ɀsv�8c�¤U�̲��ԯ��9
�@`��_��:[Ŷ�#��A�Y��g��<��ݭd��PtD��N��|�ISi���E�W�b�qU�ۜq�yf�3k�D���kwO�&뿃:�Uez�|�_.�*�fĳ�Ub9��Q�ͣZv�8�0ف��/��?���4D��l�d�y�/P(��(E�I�;�ə?�m�v�3e�������e���"M�*]3���M��u:׈S�y�է '������g�H�0͵�Fb�5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^����a$-��-C������E��"*ߛ<#
+�꘽|���]�0F�d=��0H�f�/���	%C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S�Y�8���ለ�M^�0��%�~�������˗�`�
6���.ล7[=�LAw�G�2���(��Î�HX�Iҗ��nǑ�V�3U� ��,��%r��s��B�B/"��S�Ÿ,w%��`�7.\�q�И�mJ��E|�m;ɽ�*<e�����Q��5f���$xJ���
�3"��A��ϐA��K���&Nꊓ�Hb�Tw��5�o��l �Rym�T�Iҗ��nЀ6��J���5f���>}�e�Yw*��>���>�D�'�8�����!SW��_.�*�f��vU������+C�gN��5f���$xJ���
�3"��A���q�Qy[�^N����V{c�&��N��m����������.��6d ��#��j�qKN���=��C_��K�`���/J�!#zЕ&��|JПE�[5�A��Ǽ��Yf;�b��2�w.���.�NHA�Y��g���YuI&��N���W�Xr:Z$�+�(�T	�����n��rF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�Hv@������K�}@)�v�s�ɀ&��<�o�G7�D�C󐉍��Y���%`�-�0~K���Ec�}L���R��}�Ug~	�\c�ܮ���X�%4�rY���^/�K�4�!�G8Q�d���R�Kn$Pi���!���5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�M��X�{���x,j��^̈8}�x���]L�E��uf�Oϴ���H~W�0�M1ɽ�*<e��G�����i<�R���g����v��,����
���y��Ҏ鿻�Ԡ���Vq��mK�գ�������p�L�u*�̾�~-y7�&�EO��aw��uTeR>��h�ɽ�*<e2�ڱ
�.S	����筮�>��ڻ���AoD1RMQ¥�r�֏��9��W8 �+N�����p��C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�M��X�{�����H�=L�f�5��� ����%q�qEG,��j����d�>�Mb��aO��r�Bɽ�*<e8��ꦷLX��� G�<��V�
���h���1�v,)N�	a�����p��C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�M��X�{���0{�I��X�Y6�1��6���O�>�����ɽ�*<e	��4&_)�1����G�o�O�1��q�g����������_g������� �
��� h���2��.����������ɽ�*<e2�ڱ
�&��N��O����#�LYv��,k��}����U�O4]�$ɽ�*<e*�D��|F2]�J8�F2]�J8�F2]�J8�F2]�J8�T�N�:Y�?ɽ�*<eͫ�UL��7�j8�N�d���e5��3˖>�����T����	j�֏��E��hO�99���	q����p��ɽ�*<e�<�
�F5H�r;3~��[�撴�K��֡���6���ɽ�*<eC��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�M��X�{��ɽ�*<e�n���!���D3���kf3����\�t�%ɽ�*<e �jv�5�=H�r0'�YN�`�q�g� ��1�"T4|�,�o��v���d��e�8��aڦ��ʡ7]��=�P���vz}j�笹yO$�,�ce'$��R��eL�"۠����Ks���A�@͍c�Д&b!+% �ȇj�^"�o(�E�:�::�NP��ɽ�*<e��
���ۉ�o�`�#ʓ�௝�倢���_-ɽ�*<eɽ�*<e2vr��{�l>j�m�J��}��VB�l߬�Z�Id�� �&�W���)�rc�9U�HK�ӈQQ��6P������DyMZG��K�i
��ɽ�*<e��
�����g�t��v�7��s�Z�����%��:��������ɽ�*<e�0{�I��X�Y6��a���v@)�v�J]�h���A�Y��gɽ�*<e���Ɔ��"ɽ�*<e����}cɽ�*<e1��0����,�4�+�r��y��l�VUQ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8������MP��wG��Лz���,Ȭ_@}���^ FL���0�m���ʼ��_�V�(�+ˌ�h��ܾ�uz���*��o���t��s���rĄv���0���L�
n!�<FC��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S��+�N!�W8�,�a�èr\ؾX�KX�T�����>5��Oh`	��bqI`�8U��V/� 7maH���	3Y��7 ��!Jx���]L�E�z���^B���Iy��.t���90��Z[��R¡�r��W�*�`ϭrV7��<_k�k���,(nɽ�*<e�/�����ez�,U�n[�` -A�{)����p�������I��rc嫨��~����p������,�4P�7ٝGy���FLE+����kp�l}Rk!�|F͇�*���Y�Wƍ�s(�?A�Ҏ&�Ё?m�-�,�X�Ÿ�f�2_B@�~%.DI���:��t�%2�/	J��hא�܇*9�2�\c�5��u|R���GX��a��Xڟ3�8�H�d�h���� I���}�t�wI'[]
*�J���oE����:��C�$k5p!,�7ڐ9� ��h��'i沃�Z}����Hc�9�%�\T|Aů� �B�#��t�(a�����z}�E!Ͽ���!Lؒ&�bL�.��. ����lB��,zyj���0_��A�\��B�N��%졖*��j)?��(a�����@��$�G#�ӵI�0��#Ҟ�s�-I@>������BP�\_�0'���I"ʈ�W�rB�������i0aXK��2��H����D���i�6 ��Z�)a��\ `L���c��}W�R�#C,��n�Yx���|��/_��P��r�k���g��� H]K�s��K���{T��
�7`�	�6�#'	��m�:��eH��J�	��[W�DC�"�N�?�ot�'��#~D��\��KB����VL��'�s���7K�f*���b�0qK�s��D�1d�	!4wI�o P��z9����D�����e�mu���H��H�
:��p��؋9i�^��,1DԾ����\J���H�.'a:�s�c�A �Ы���VI#�1z���x�q��Ǝ�b\[��½�#��$̆���5��0^v�'-�r�D��6�^i~��b!�t�&��9W����z��\(u���?�9�o<̀�t����{����f�2_B@�~%.DI���:��t�%2�/	J��hא�܇r���+9}�t����{����f�2_B@:P��dS	nT��e�&��F]�J�������	U�֝�%��LP�b�I�hS\'��/���`b]P�L��ϰ�9_��]-͍)�,\���� I���X�%���=��dn'y&̢���N���ꗳ�)�7��y���#H����^'�2����:W�0s�����S�_>gN�-�:'��$+���G(����^Le�0�[��z����jcbb_�B�,��y8f���B6Km���'�5uEq_�<|7.���|N;X�^�I�[\o|�o�����|"ÝW}�utiO����+�%�Q)=d���E@�׺�F�b3��5����4�fgHg)%�RPz
2����$_�>U�V-'�I��.3	
.5�4w���
ק5�C>��M ˶�{T��
�7`�	�6�#'	��m�:��eH��J�	��[W�DC�"�N�?�ot�'��#~D��\��KB����VL��'�s���7K�f*���b�0qK�s��D�1d�	!4wI�o P��z9����D�����e�mu���H��H�
:��p��؋9i��������a:�#�f"�6]v��P��w�	|"�@Ҍp���O��"P)�6�m�`�� P����Y6Z����*y����,��/�&�5K}�*���ՙ��e'�������s�SŠ��z��Qd_No���?�%6=�N����:��*D�)�=��x�Ϟep�h0����p��a!�atXCB?�<X�aҥ���4f<W��ג$OJ�7� ���7`�&5��=��od2p[�������Ɯ�h��e��9ʡ�όT(ɇ�qkaDt¨���:!�6AD6B�iٲc�z��+��+T��L��l�����O�l�[#�e�F2]�J8�F2]�J8�F2]�J8�F2]�J8�]^�h����T�rD�G�9#�xS��*�N�S���"l�c�"��%�mƚ����vW�,Fu���Hl���͆��7�Z<e����mAd[30��4!�6�?����2�^b�����a�DQ�BE�?�Ҥ�a� g &��m �w�3��4��?#|{��i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8��"�iS{/E�́7�׈�|�.�Q>���ě�T�t�g����i{WU��q�����b��i��<�a�]���-�几��p~rևzϯ=yu����1����bT�>��*�����j���R#l��凉�k����_P!_�V�����Hw^���]������˺����i$�BMo�A�T� �{*o��^��DF��t)vD�厜1g']5��kL���RI?�st��}~�M,�Q�.#��W*͓M�7@^|8�f��j^�C �<�CB�\�u�<T_2��G�= D��VZF��m����9�@���1���?�~ �(	o��P������d[�� �=�;���*����t=X��Q�k��/�����V��U?��4�&,䖼��X�*f��p~rև}��~�����@��W��Q��t$�����%�R#l��凉�k����_P!_O�4�WW�hHw^���]������˺����i$�BMo-�lI~�{*o��^��DF��t)vD�厜1g']5��kL���RI?��@ۃ��\�u�<T_2��G�= D��VZF��m��C\!���X��t=X��Q�k��/�����V��U?��4�� �W���������%�R#l��凉�k����_P!_(�a"£� {*o��^��DF��t)vD�厜1g']5��kL���RI?�5~�tC��!\�u�<T_2��G�= D��VZF��m��Q�-/����t=X��Q�k��/� P���t�	+�V��m��SS{���r���4GHd��>!H7���.%�R#l��dJ<R�[��68�Fxɽ�*<eɽ�*<e�V�w��~]�������v�2K� i�� �=�;���W��5Y�ɽ�*<e{*o��^��DF��t1�n��gEaTq�A�i�b�=7|�ɽ�*<eW��_��_M,�Q�.#��_.�*L�#�I~�#鳼F
�sf8~�^+����~?MA��1���?�~ h�z�3E�i$�BMo��u�MЌ��aRI )��������t=X��Q�k��/�Gf���<���_P!_ҍ���I]��~^-C|��v�&�����F2]�J8�F2]�J8�F2]�J8�F2]�J8��� �z F71��!{B�)HA�+��^큷����X�vI9���	��3I��N�^�5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8��B/P �S�Ͳ�����v��l�P��yl2���f��S��<l���P�]�9i�eE�P_��1�]�Ҽ�w	�x�Ae�+Ss���Y�|���~��WfAϟ�o�	ɘoƩ��-I��a�����!ܶ�5��Oh`�}G �}���E϶1w��%�mƚ����j0��;�"�����Ͳ�������0%�[�yl2���f��S��<ٚn0��.>]�9i�eE�����*�"�����Ͳ����d�(���c5��Oh`�}G �}��&H���^��~��WfAϟ�o�	�>�CM k]�9i�eEѢ�yO��"�����Ͳ�����ƿC+��5��Oh`�}G �}����q46�e]�Ҽ�w	�x�Ae�+S.	o�L���"�����Ͳ�����cI�u�0��,�A�#-I��a��s�Z�7z�A�IlHL]�9i�eE��d4�fl���w:3�|�%�mƚ��p�>u�b��/�+d����~��W�����O�i��S�yl2���\��b�|��������5��Oh`�}G �}�,�K� ^]�Ҽ�w	�x�Ae�+SpF�3�[9~�"�����Ͳ�����cI�u�0Ǫh5��P�]�9i�eE��d4�fl�ne�� �m��~��W����h=$"<i5��Oh`�}G �}�٩���Ò�"�����Ͳ�����cI�u�0�����a��]�9i�eE��d4�flǇ������5��Oh`+�Ct��0�ic��ݤ���b���\�V'Ba6j�؋$��,!����9��\��b�|���?���a���z��I��#U#*�[�jtKϒwfյ�J���.���w�&�u��;�����A\�7�nr�����g�Ә����n�F�J�ʛm_���r���PY����*�U���	���vq�s3����n0��?�i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8��AP~�;����I��AG#�x��v��}g<A�:�X]��V�X�˄���<��q��q8I�x+qjy|�'��Y�n�K�m����F�rJ���C���}X�1�{��F2]�J8�F2]�J8�F2]�J8�~�&T�S�=c@�LT�O�W��̴%[�{���`��6Uw��JYw�8�r�rz��ښ�Fȧ8����צ ��Q�E�]f�1�m2\,�����g']5��kLDQǺ��@ys�w\6kznr������G�t:�~,��ՙK���3'L�S'��������}�y� a�TaS�W�k�}��(p���i$�BMo�����dAt��I��3N����v4�����n�*��IYk��S�1O������R�J���}�0״���y�\�i��<w�W#�+X�$�rҞ��Ri���	7\��ہɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e����6wFlJ@Ҷ#�hMU)�_>$'��PSɽ�*<eɽ�*<eɽ�*<eɽ�*<e�/���%�����p��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�m�F�(lJ@Ҷ#�hMU)�_>�Ri����	�nɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e������a>�;5_s1�E(�p&�~^i�ɪ*xjaL�	��:��=X�-��l�!v.�� ����3ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e����6wFlJ@Ҷ#�hMU)�_>l������_y� a�TaS�W�k�}�I ���ؓi$�BMo�����dA�F�N��J�	x>��/����C��Tɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e`������Zݪ+i(�'h(����+NII���F���b�i$�BMo��u�MЌ��aRI 	q�ho?�����F2]�J8�F2]�J8�F2]�J8�F2]�J8��
�%T��sx�6F�`��Ut'����('�=�3����^����W���[�&,��z�r@��YH1V'Ba6j���u�ԏU�H���4��d4�fl��8����iͶe������*��J����9 �K��m'WM��>n�
���lį�X{�g��K6��+�?��0���]�ͮ9�!����cMOd���.����p$.���km]sQ7Oq(�b�ٍ�W �-�] h��^��}C��v��ɽ�*<e=Hg�i�|C���P�s���bg���{v���ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�1��$����7��_��*���m��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�]D��ˁ�s�
��-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^�M��?��it�am@
��&��ͳ��};��=��c-X�-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^}��Pj���e"����s��N���c^C��ɽ�*<eɽ�*<eɽ�*<eR��z��#A����k�ɽ�*<eɽ�*<eɽ�*<e��_��l�A�,��p���Yr5ɽ�*<eɽ�*<eɽ�*<efAϟ�o�	6�����aɽ�*<eɽ�*<eɽ�*<e`ύ���#Si:� ��Bɽ�*<eɽ�*<eɽ�*<e�i{ޝ��i�B:�F�d)6�!��ɽ�*<eɽ�*<eɽ�*<ef��S��<�@�a��5ɽ�*<eɽ�*<eɽ�*<e7��� h��U>��[{����p��ɽ�*<eɽ�*<evS+ё@��j0��;����_��ɽ�*<eɽ�*<eɽ�*<eR��z��#�M��$�,ɽ�*<eɽ�*<eɽ�*<e��_��l�-��k���Yr5ɽ�*<eɽ�*<eɽ�*<efAϟ�o�	G��$�f�Mɽ�*<eɽ�*<eɽ�*<e7��� h[}Y�����Yr5ɽ�*<eɽ�*<eɽ�*<efAϟ�o�	�����\Zsɽ�*<eɽ�*<eɽ�*<e7��� h�HdE�����Yr5ɽ�*<eɽ�*<eɽ�*<efAϟ�o�	x� �Ͷ�ɽ�*<eɽ�*<eɽ�*<e7��� hn3�Ė��ɽ�*<eɽ�*<eɽ�*<eY�5��y�)�����Q��c���-p�>u�b���?c���ɽ�*<eɽ�*<eɽ�*<e�u_�2�P}�ko���@��W��ӆ�uN�)�*8rB��p�>u�b��L/`�Z+�tFK��Xɽ�*<eɽ�*<eɽ�*<e�u_�2�P}�ko���@��W�g���Ǭ���*8rB��p�>u�b��{�\t�O+�tFK��Xɽ�*<eɽ�*<eɽ�*<e�u_�2�P}�ko���@��W�R%Љ_����*8rB��p�>u�b�58����b+�tFK��Xɽ�*<eɽ�*<eɽ�*<e�u_�2�P}�ko���@��W�ǗH4�g%�*8rB��p�>u�b����R���+�tFK��Xɽ�*<eɽ�*<eɽ�*<e�u_�2�P}�ko���@��W����?D���*8rB��p�>u�b���Y�`
�+�tFK��Xɽ�*<eɽ�*<eɽ�*<e�u_�2�P}�ko���@��W�Ǹ���]�*8rB��p�>u�b�ܴ��95+�tFK��Xɽ�*<eɽ�*<eɽ�*<e�u_�2�P}�ko���@��W�q����'��*8rB��p�>u�b�Cyڻ��+�tFK��Xɽ�*<eɽ�*<eɽ�*<e�u_�2�P}�ko���@��W��Q��t$�*8rB��p�>u�b�U��z��+�tFK��Xɽ�*<eɽ�*<eɽ�*<e�u_�2�P}�ko���@��W�/�{��r��*8rB��p�>u�b��%����+�tFK��Xɽ�*<eɽ�*<eɽ�*<e�u_�2�P}�ko���@��W���TS���*8rB��p�>u�b�U��E��+�tFK��Xɽ�*<eɽ�*<eɽ�*<e�u_�2�P}�ko���@��W��+	0�
a�X��f�����JMWs��+�hh�@��|v�|�ɽ�*<eɽ�*<eɽ�*<e�GY�fX&�i$�BMo�A�T� ��M~�7���a���ym��Z�1��^��H�Ȣ�������*ɽ�*<eɽ�*<eɽ�*<e���}��$�7@^|8�f��j^�C	%8���v0�p����cI�u�04D��b$�a��[��ɽ�*<eɽ�*<eɽ�*<e����%������d[�� �=�;�Ա3��.N6�He�����d4�fl��= �9�+�tFK��Xɽ�*<eɽ�*<eɽ�*<e�u_�2�P}�ko���@��W����(�F;ȗX��f��������g|��+�hh�@��|v�|�ɽ�*<eɽ�*<eɽ�*<e�GY�fX&�i$�BMo�A�T� ��@N���?�a���ym.�^�<�e^��H�Ȣ��Yr5ɽ�*<eɽ�*<e��I�v�:�>&��l-�i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�YZ͆ˎ������!8t>�y���_�ޔ�~M/*�t��j��|9����@AVKyO�\13̭i.�-�"�Ac�;7�k���C���*�zðɆ��q&�:=�-���G)�6� Ri�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8��ob���O���-��ѳ1<�+͓LBϏ�ݸ���RE�C��&���	B�9��U��@g']5��kLvA���8E�0{�U������'��ߔG�=��}��Pj�s`Bs	Nx>��4�3�\���e"���|{5���kwO�&뿃�5��X���d4�fl�\�`pWvcT	����as�Z�7z࡟qn8��?��<��ݭ.苢��w�ɽ�*<e�{M��?��~�B�ʇ��t�i|�����N���Q�)y����p�����f���:ɽ�*<e�K��r�����n�y��;������cW�,��Wz��rkά�
è��$�;Wd� �=�;���W��5Y�c� �a>������YD��Q��e��"4�R��׾ɽ�*<e����j��{�.��]����p���
��2ˀF+�n�/�G���Xv�kջY@f����cW��H��g澅���Ȇ�'b1A�/���lco8����cW��H��g�V'Ba6j��se�gې�d����pھi��͗
U�H���jp���{���Ҥ�b�~��r�Y�(�&�o��� Cb=��K�X�$��-5B�f��<j9D�m��j��_h�-?�68�Fx���o��c/���Y�Gɽ�*<e�O5l�u`�xK���6{��I�u"�#���{���j?�%BN[VL�
D�2���2S'L����%nP��cɽ�*<e�.&ׯ��1? ��6�5���@Ԁɽ�*<e�<�DR��ܞ@/��`nQ���-x�cI�u�0���V�uCM+�n�/�G���N.�b���ya\Dà��������3٥���p�Yf�{��t��;��f#Y���LT`�(O��y�~�k��v����7l���@��W����<,�,{H
ʢd�ԟO���<���I�h�K� �=�;��nO���ɽ�*<eɽ�*<e���
����I�h�K� �=�;��ڽ�R!&��y��Y�ޖ��r���PY����*�UԘړ#4^XE�s3����Qz^�j~kk���,(n���h3���*�Ӈ�k���,(nɽ�*<e���N.�bs���!�1U�PiD�VC_��޶(:vS+ё@p�>u�b�p"�opO���O���WA�Y��g����,�4r�֏��9�&TO��A��%���]B]�-p8�?��שePY�$s-�E���dx�$�i$�BMo�}n(Y��x{����ߔG�=����YH1V'Ba6j����<O_ɽ�*<e�{M��?��~�B�ʇ��t�i|�����N���Q�)y����p�����f���:ɽ�*<e�K��r�����n�y2H�u� ^�p���ɽ�*<e���gR��8Uc1/�ɽ�*<eھi��͗
nM8��?�4�pK�ݦ�k�ļ�*���%nP��cɽ�*<e�.&ׯ��1? ��6�5���@Ԁɽ�*<e�<�DR��|d�fO~bA�!\e���(rd3��ɽ�*<e��;?Q3Ց �D:X�m�׻\-�!���s��U���I�v�:�ߔG�=��'4M���/v`S^!������·i{ޝ��i�!]�?T�Rkc��*2�r���Y���A�Y��g�i{ޝ��i��V�X�˄kc��*2�rX 0),�xn����p�����Ɔ��"����,�4�����n��XS�<)�	~`v��YT	������z�V���p�(�bR0-����!�Np�>u��9������/�žC��Q�:�`�&5�^��_�ϻ�u#_��I��_?�w�G��7�H�+��	�R�ܛɧ4��pJ�rC�hbP�7ٝGy����d��X����G���R�ʹXr�G�Uk���x���]L�E�؝�Bb�a���o{
��~�H��V�ԛQ�Kuש���q���e��QRp�5�!�b�a�¸q3:ɽ�*<e!Bÿ�L�������
?�	�Ù	�^V̷��Ż=͈�S��eH���Ù��Գ���P�s`Bs	Nx��M'���V�6���f�I4�������9A�Klײ��:�#�y����o�:���:P�,���QI�`V�f�BvS+ё@�! ���9����5��e�t���>ٍ�W �-�] h��^���QCYlþoD��[�_o��u�삙��q�E������b"���	t�nQ�ɽ�*<e�*�GP��tXCB?�<���A�53�m~�ƪ�J����a-��}�N;�ԉB�'╆G�Xz�(�Ց5�^V��&�������p��v�ُ��HS�Mh�7^qYj��gǧ��3P)3�����
C�ܤɢ�]A.�I��oQN�ɖY׎�Һ��F�Y�zU@�iL�k���,(n=Hg�i�|C���P����{��s�V��n�T(��! ���9ƪ�J����&r��/?��� ���U[�ԩ�Q���������,�4�
�9����W}��Z�5�1�`Ӧ�g�'*
��� �/�OՖN�~)�X��޸,�Zu�;��)�#[�:Q��"7g��衅��:_���5��6��u*XdE�z6}ȭ��5&��#fH����=<�K8#��'+dL�9�N��|Uw6a���������"Uy��\�V�W�v#@Y�����\��&�������p��H4���{M��?��~�B�ʇ��t�i��H�Z�2�r�\L�sR#���	T�9���8�a�bzHٜ��IA�l�%!I=W���A�>�l-��ɽ�*<e�0Fct���H�M��hI�t������<��GoT������WE��@��ɽ�*<e�$�i��n�}\��'�}��9��\!����ɽ�*<e䧓� 2��.?�$R��&�/ n�^5)��ɽ�*<ed`�.�Zyar�}��׭�7��_���H
E#LPA�Y��g�������w��Sk�jQ!I=W�����t���U����n�fɽ�*<e_���#�*c�H�M��hI�t�������-�8wɽ�*<e��=Lc�H0�J:�3WQQ�g��.2P:���[����p��n��c��=���<�! ���9�.�>Ƒ��d񱔟�A�0>��2ɽ�*<eW�VegW����7!#�WQQ�g��.2P:���[����p�������9��ߔG�=��@�^�~=����(yy��*��o��L�&D��7��_���n�3�81��i$�BMo�D˟]e�zN϶ήh5��jqA��|���Ũ7lɽ�*<eJ�.4��X��]D��ˁ�Er�L��<��GoT������WE��@��ɽ�*<e���И��S�k:�Q�"}��9�&���[-;��G� �Ԭc%�ل��pľ��ɽ�*<e !g�T�]D��ˁ�Er�L��<��GoTO�s�滛� �/�OՖ�;�]����zb|pm���x�z��\�J�$��kF`!�@,�Xڟ3�8����!��<,�Ŋ�5�+��:S��؜!��'����t���UY�/�YP{��s���pľ��ɽ�*<e�k�\�!�g��#+��̝Er�L����-�8w'$��R��e��Ω-b��v��,�����h3���*�Ӈ�k���,(n7��� h�p��q��!I=W��ɏI6�� &G7��� h ��O�ט����dRݒy~O�5��5���Ɔ��"����,�4����/ַ0���(��A��mt�[� ܢ�:{��yO]�&��I���R��A|`�$������kȡ�B,ŭ_
j�����ͬT$OeMS���s�C�罤�9.�f�i����
D��H7����{�ƥUuh��V�g5D�l��9q�X�:׮�5:��KL����z�>�4[���{u�^ק��}�{�ʘ��SD!��Ю���0�V�٦�����2���X�����wD`֡��y����"�m���F^��`���#H����^'�2����:W�0s�����S�_>gN�-�:'��$+���G(����^Le�0�[��z����jcbb_�B�,��y8f���B6Km���'�5uEq_�<|7.���|N;X�^�I�[\o|�o�����|"ÝW}�utiO����+�%�Q)=d���E,��h��DZ�x���F\��w�0��8w���c�Y�l�%�tB�*��� �&&s�:v3�9?k����Q������L�����p�N_�qe�
��>̊��%�
�T���k���g���*�F/��q+�\��$|?G��a�G�x�D�9ϑm�eQ���9*Q����� P�7+��$-���G[�z�A��ie�\#�_Hc����'d����uC)�E���Q�0)Dm*
kma��ݑ�`��N��X5/�)I�|��o9�H[��UF�n]h�^�o��p����=����+P
���(�5;B�W��M��v��E�`�w$�P��j�:�mheˣ��:��?Dg,2ms����{Ue#Ty� �I�quȯ����2���Ե+�ynB�;{�7�$$x<nҤ�b�~��Mg�������#yc{]�ͻlU����\�IFa���o{
��~��i��܁�q f�&�2=�&�ظ���tk���}Ո�,�AQ]�h�j�v���� ��B迅9DԄ�r7uo)V�&�>\���^��0*eL���J:Գ�5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��x�7��ʎJx��{昁�.��Jm�X���F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��
�[o��=�	rr���6�XoN��5+}4���5�}�'�`�&5�^��_�όB��N5��8B`}�wG��L�qM,�Q�.#��Z�j��xK����M+DW����DF��t�.^)C�q*L	��D2h�n�3�5��Oh`o�s�Ъ-��ڽ)n���V�²z<r������" �ΜH9c���0��hf�%��}�F/�zo��&�{NcB����J:]_ʈ��k�y����<o��s�Xq��hH��eF9YH,���N.�b�k�h��C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q��"
�F��^���.�֋�
�j: S|s]7f�q9�	��6m8�W8�×,3a[�mf���~;�_@���ʇ��t�i8��x�z�d�H�Z��9B�ˎ�U�|6f�aA��n3����p�n�`U/�G<Ih.��<��� �{0˵s����)t\��?�n�1Rb �v!�(��UO���.������V���r)bgdW�yz-�՜�I@j�ZC��Ib[�഑���'~q��s�s%�=4RӁf��Q��|b��g��[B����W�B�*!�nUrW��_s2j9�gi�Vo�Á�\ gS�!�ex��{m�tst�������r;m ��H�$r(�ÎVnZ����u���	�P�2Sn섮�rS��������C�?�򯁣��A��4y&G�-��W���޵7C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q�݊[ĩJ2�\SG6��T�*�����L��&�e�S$Ҥ�b�~��r�Y�(�&�o��� C��o18����ؖ�8��ŏ>���b`�&5�^��_�ϻ�u#_��I����?"q�	�&��Xƻ�2��{�׻poH�����20rY�1���o�ߔG�=��C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q������n��rT��M���^��_��C[&0q����r����y^��_��zd���VJUT���i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��l��q�'4M���//�%
q�sڝ�o� }�uKO��m2�6]�9����Y���k����� �
����+(M�e~���Y���k������ɽ�*<eQ3��Ѓ������
?�	�Ù	�^VqYj��g�K�����J�rC�hbɽ�*<eɽ�*<e�{M��?��~�B�ʇ��t�i��H�Z�J^o���.2P:���[����p����8t������p���_F��x�J��E|�m;ɽ�*<eɽ�*<e�{M��?��~�B�ʇ��t�i��H�Z"��i�?Y���:����|�}��������
?�	�Ù	�^V~Z��~��)�T��ut�hA�Y��gɽ�*<eQ3��Ѓ������
?�	�Ù	�^V~Z��~��)�1dW�*����g���ɽ�*<e�؝�Bb�a���o{
��~�H��V�ԛQ�Kuש��t�V�,��{M��?��~�B�ʇ��t�i��H�Z�=���߿pɽ�*<eP�7ٝGy�ɽ�*<e9�ݞR��=�j�8]����Ĭp{��p��q���{M��?��~�B�ʇ��t�i��H�Z/�I�|����O��ErG�Y�tѥE��䅓�g [pe�2�f?*�D��|F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^,4���?w��yj��oy^��_��C[&0q����r����y^��_��zd���VJUT���i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��l��q�'4M���//�%
q�s���]�[�JПE�[5ɽ�*<eQ3��Ѓ������
?�	�Ù	�^V~Z��~��)�O!��##��$�ŹCktXCB?�<���A�53�m~�ƪ�J����K�O!�V,\�$V �0�ɽ�*<e�{M��?��~�B�ʇ��t�i��H�Z"��i�?,Y�F���fAϟ�o�	A�Y��g���{���Ҥ�b�~��r�Y�(�&�o��� C��o18��x�J�=bX_�T�t�g����i3� (qɆ��q&�:����\��ȷ���Q�����p�����Ɔ��"(��Î�HXo� T�uїJ��\��Jx�T�t�g����i3� (qɆ��q&�:����\���&�ٵ{����1��0Q���'�}�qTeM���=E��Rx��w1X���yO]�&��I���R��A|`�$������kȡ�B,ŭ_
j�����ͬT$OeMS���s�C�罤�9.�f�i����
D��H7����{�ƥUuh��V�g5D�l��9q�X�:׮�5:��KL����z�>�4[���{u�^ק��}�{�ʘ��SD!��Ю���0�V�٦�����2���X�����wD`֡��y����"�m���F^��`���#H����^'�2����:W�0s�����S�_>gN�-�:'��$+���G(����^Le�0�[��z����jcbb_�B�,��y8f���B6Km���'�5uEq_�<|7.���|N;X�^�I�[\o|�o�����|"ÝW}�utiO����+�%�Q)=d���E,��h��DZ�x���F\��w�0��8w���c�Y�l�%�tB�*��� �&&s�:v3�9?k����Q������L�����p�N_�qe�
��>̊��%�
�T���k���g���*�F/��q+�\��$|?G��a�G�x�D�9ϑm�eQ���9*Q����� P�7+��$-���G[�z�A��ie�\#�_Hc����'d����uC)�E���Q�0)Dm*
kma��ݑ�`��N��X5/�)I�|��o9�H[��UF�n]h�^�o��p����=����+P
���(�5;B�W��M��v��E�`�w$�P��j�:�mheˣ��:��?Dg,2ms����{Ue#Ty� �I�quȯ����2��ȿ���&�C�16�wX �V'G��>E7��`��3�����h�O1>�BɆ��q&�:	�5zh�O1>�BɆ��q&�:�O�|Bۡ�x�*B��0�ѡlv����լ-:��I���v�`E�bΨ�c�꺉�@jB��Z�!��3Sr1�p��*��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8���g�7y��.�NCE��A�ώ1�Đ���A�P��ĬjCˬ�eQ�cג$OJ�7�,�w�͉�%)��f8�X��"u)mT.��AVKyO�\1N�,�9�*�F��+��Ɇ��q&�:�P��]��Zg(~��Id������ɽ�*<ei'~���ѯ2ZF���f^��_�ϕ$u�;X�."aJyl�� ?�}�سodI%C���0Q�.�?�(<���l-�ɋ�;�n�����Д���DІǦ/FO�u&7/��b��F��ޓυ������^f?�(<���\c��tҤ(��7���~yڛ��P��Y+z@��tCp�h6%
(��<����L������:j���+��!$k�3M�(D�n�<�?�(<�����z�џեAB��d�x����2+�j����S�>+��	z���J���a4�a��>�����i͆:8
'�J�r�E���#v˂�Wi��p��"6%��n���x��p\g�2�m�<�7:��@P�?�(<��Ҩ� E�k"����Z���X!9KҮ
��q������C�Jl��xhϱ�ж�Ⱥ�?�(<��{��~���8U+q��<,�gS���h������+��Rpv����@OQr�ɽ�*<e�Qӑ�y��Ebk�&�8U+q��<,�gS���h��r��c�{��Men:5�ɽ�*<e�X����l`��{�`t��MG9�	�(kC;�,O�]�o��@ ��'��;<��݋�ɽ�*<ex��8 �R�nq��q\B��;Jq�S���[���`C;ig��XWaMڶ������옙9�W�\O#AY�s)B�?1�4��ߤ^�N3�"d�D�`(}QM�Eiv/d��dK�����N�����_��d���t�Q}���-����m\Ʒsa
���������b!TN������*W�=�oE�V��1��m$�aܔ�H$mK�{B�a�!n�y��G�[ �&��������*|&حF�ù=#.|�C�� d��5�v��`p�U��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�4)�}Uh���"ﾆ��78	�*ޮ/�8�:o��
[z�Ţ-���f�o��� Cbv�A:C�]�ͻlU��]@x0�z�ɽ�*<eɽ�*<eɽ�*<e:j���+��5=d~5�ɽ�*<eɽ�*<eɽ�*<e��_��l�ȸMzvwɽ�*<eɽ�*<eɽ�*<e�E�a�*SB�:وR��ɽ�*<eɽ�*<eɽ�*<eK�Bѫ3�0��N��~ɽ�*<eɽ�*<eɽ�*<eU�H���jp]�������������L��ڞj��J'�bPw�<��'���Ι��;%j�q��:7��Q�k��/ޏ����[@�.�1�7Sa�.U�[�x�����i(��ï�V�E�y� ������2<�j�JW����iR~�	4�դ ����E�괓O��d���5����)@��v,� +��><�Ҧ �l�CЉ:�I�/�Yik�}$xS�"�]),Q���p��S=�~���]}���C���-�u4��[k�H|@������[rhY[v�_�>d�Lvl��\|��c�q%Wr+�1<m#�:�������O��y^��_���5@xɦ\V��L�̨˼h:�?a t�oe0vZ��v�hN��W�B�����B� NM{9q�����R!�	{�b;�^:S(��g�}	}@�PrR�v��8\����.i �e�z�,LM\��S�F��êT �ʇ��t�i����G��ɽ�*<epa�{P��er"�|��&�|?:g�E<��(�|�wk����3爸��I�Rl����4\��&�QÀnG�:4N�₏����s{��O�FnE];hi!�����4���d����uT�ڞW�A��XW0��/��acf�b%���z��8EWG��sAd���l/@N�~Nd!~5ꦋ��C�_d���""9���z��R�K��:�>S?�����.����REi� SO�r���#����/b�r�m0{���"���ޫyw���2vl�n�h��+_���Y�.�)��lk�a$ejˑ���W'�d���p%(�,�Du/ndZ���ruČ�!�҄��;$睖�� U�0;���m�IτM=��:⍁��6HfiF�JA��G��.s�x�ZG?��6���BrW��mVW��c�=�����[���!�Np�>�`V�f�BO�
�����̻U�QHi�Yex�����p��O��B!BX�`8gim�ڔ8GR�
?�	��9
�/��(��)��ش8��L�-���M��o H�'���8t��0.d�չ�R�f.��d��Z���9��_�ޔ�~Mفc�Qp�yq�(����'�i����
��j�,�1������b�H�A/���*Hⵁ����@��\�l]��G��犓I���$+���G(�bg�y��#A<TuX]�<r�k������9�,ޤ�>�����3vB@#���R���׉:ƄkC<�mo������<#�<{M��Uh�Y�h���Oܗ�q��	~�������-�p��"y�
5��	x>��/��zg�b%�զe�R��I�f���W�h83�fJ#j�S������vE�����wm~�������^	+��Т�M����с-���N�ʆQ'�m��=3�E�w�z��p��u��d���+ԓN��6�Wȵ�xf��TP��7ή�Q%�!��6��6�zKhl��R�]$b�-�@� �!feY�WȚ�j�hx���]L�E��]{X���Y�V'�P���=����{:���+�fOKPl&�,m�E���p�9���Q�D�[r�P����n�L�P�`�}9���^��TfzFj`▘9�����V���rzM=��`V�f�BO�
�����p��V�e�><��P%vS+ё@	���!R��RW��OD	��݊��T���#�X�7�_F��x�gƧ)������7cO&(Pط�*EMߛ'!���9�ݞR��=��Ic`�JN������ DO�򮾋.q�-��-�5�e@�Yk�Wx��Z؄Tڴz�6|"��K����G���R�ʹXr�I,N��o+m��Fo�lS_O��k���,(n3ƹq�nNso~����&�p�'��7��E�a�*S(|9���XI��9��ܰ��7���G��m��	L!�v�7A�Y��gzu�V�����E�a�*S(|9���XIˍ��V�!�v��,��j`▘9�����VA�/�l<~O~���h�M͠8�H`�����o���������U�8�s]�����gL�y�q�!�g��x���h�H$t�����[@��ny��_������
:��{g�_F��x�gƧ)������׺uB*��-�^��{p�� GN��%���K��`��r�@��ӂ�7����I��cW�n2dꜱ+�	���k˽".$�WFi�U}���7��&�]���j`▘9�����VA�/�l<~O~���h�M͠8�H`�����o��������O�
�����p��V�e2F�j3ɽ�*<e�g��x����*�om[t���y�Pɽ�*<eC-����ɽ�*<eq!yt���ZVt������p��3��֪��	D�ܣ{U]	ȳ�ؾ�k2�G�Cz\�@bn���=r?�eƵ��&�㥷��{��߂]0;�G�	�M��)��3�uѨ�<��!����;��pY$x���]L�Eɽ�*<eݕGء���`T��4�@r���28ɽ�*<eyW.�Mˎ��O�pٺe�ɽ�*<eAN$(��5ɽ�*<e�g��x��Ċ�7�tvTa�upIf�{��t�����/ַw��g�.S�l�Z��&��!*�,;E��O��]�Q}/��<��P>8X�QX�ck�X2g����Q�e��!���x�[Pm��wr�]�e>��p�!���bP�"Uy��\��P��{þ�/�žC���U�8�s5l�UK���4[|���@��X�xhp0��ᏺ�z�y!-x�z�����'ck���,(n;N{/�~:|��`@�&Q~�0�n�����|J&j��m\Ʒsa
��������bU�Tz����ǁ�T���|\d+7�s�O(~�Աz�:��0�*I�p���b�!כ+�r��y�h{O�v;��eg�@��d��J^��Ҧ �l�CЀ_�`��'��-<���AIVk�'r-ײ��d�����ANφqy쎤d�w�r����r�j<ڪ��Ca�֥�Ѭ:�W]��Z}TG���������0��O�&Y��_�:��+��k2�G�Cz\�@bn���=r?�e�><��P%O�
�����̻U�Qg
��V������j`▘9�����VA�/�l<~O~���h�M͠8�H`�����o������� �
����+(M�e~����d�L�����p���E�a�*S9W��)!rِ�M�p8�b3,�i
$�ɽ�*<e�.U�[�x�ɽ�*<eC-����ɽ�*<e�)��8t�d���t�:_C
�V[�T��%z�ɽ�*<e�&Nꊓ�HL�"۠��JПE�[5kwO�&뿃"�9u��夣�P1޸��ϝ<��Uצt��y4��"���JПE�[5ɽ�*<e���M���Nl1p�N6&�9_��Rɽ�*<e�)��8t�d��t���I�2�9��`1y��V�7Uɽ�*<eC-����ɽ�*<e�)��8t�d��3`�P�2�1,���ʽ���⼲��;�
'$��R��e�����kV��+�r��y�Q���'�}� �M�Y�8�����Cz��(I�����[@�?���|��
���M����4��Is8��/�žC���h3��.
�_F��D��k��-�]d���)%��b0�δ�C:Z���/�žC����@�������N�	��FMg���Yr5ɽ�*<e}�>�4)=P�eP�H.�I��oQNɽ�*<eG��.s�xɽ�*<ezu�V����ɽ�*<e��h��l� �0�9h��)τN5�G���8t��ɽ�*<e��Yr5��<��ݭ�`V�f�Bɽ�*<e����q�E���蟣��B�3/�.��+�>���1AiD�`V�f�Bɽ�*<e3ƹq�nNso~����&�p�'��7�ɽ�*<e��h��l��G�i�O�;t��5�92�w@����;kɽ�*<ezu�V����ɽ�*<e��h��l���kO��~&������vxϕ�o��â>"@�ɽ�*<e1��0����,�4����0b��*��-`������Q��5��9��O�<B��u �?Pƅ�i�MNkT��ߡp�㙞ɽ�*<eɽ�*<e�J4�2�|�� HA�M�5x�R�F�hԚԾ3�81R�c���2p[�������Ɯ�he�[�Q��$x�"������^�_<��e�u4g��2ޔ��Vn�{#��I=��cП�%���[[����%�#p����?�[�#a6駹U������2���Tu s�_f9��1���nxr�^���Z�a�Es�������?_Gߨ,��4c7���˦U�5c(W�-� h�����\zӄ�Y������t���,Y�^e[��z��I-듈�<�����שG�P���8B`}�FW,P���O�B�]t�Jg����ͮ��&T�A�vb!��wF�Q�k��/�a),5�,z2�n
2�r)f�h�P�m�p~rև��}G�5�X�%C���W球&�� �ϵ%[��zN�����M7@dN� 8
�Yۺɽ�*<eҝ[��R���r�<xAY{�#w�)3��Z������@d�����4�)�_π�;�A�-� �z+\�`둺��r�H9�����Җ LF�6ҷ�׸�3�q�w��ݹE�=5�4��^��l�ҝ[��R�� �3Y�S��%�>v;�e�`䷟����{v���j�������	�;�;��H3�=�Xx�\�uɽ�*<e��]/߷�WW���;��X z_.?�PZ�����ń� �3Y�Sl�7ñz�ɽ�*<e�����+�n�/�G�w3<� j z_.?�PZ�����ń� �3Y�S��Y����ɽ�*<e�����+�n�/�Gl� �J�����Җ LF�6ҷ�׸�3�q�w���LQ{D���8��8ҝ[��R�ɽ�*<e�4ł���#OˬzO�I�D�J�ɽ�*<ei�OϿY�M�L>�;>c���D%��ɽ�*<eZi��LύE��9��h.g�/�B�VT�́8�1���E�i��\;�&��z�IYLy'�~#��ɽ�*<e���U�&4��%e�܉X�X���H{T�_0��ݑ����V_^��k)ɬ׼W��#T�q��H�ݐ�ɽ�*<eY�I����b\	y`��V�mB���x��{}�����;��ɵF1���*l����⃦�q��i��\;�&�[.�[���uZ1��������ZEŝ�h8=�d&t$���9䌒��A�B�dl��R���7R��M�m��H� 3�`?,D�}ߓgߙM�9gul�@2��+��c��-F<�!����?�JϽy��W�h��b���csu�GA����mr�B�j��O\��v������y���5_m�������w�$=�d&t$���9䌒��A�B򜈱���рE������-F<�!����?�J\e񧏟5�����Z_O�gOO��Ctb %+�>|
ϒ��޴W�����ɽ�*<eɽ�*<e���B��n��W��2���m���_B}���M`.�m`�| ���O�QMyO����u���2nq�Ř�x`һaB�ɽ�*<eɽ�*<eGAȖH1����!܎^R��l�G�䗋��[0����E'bwE�m`�| �fN��ʷrP����u����Q(�>·�ۃRIɽ�*<eɽ�*<e	�9
G���[4@���}6�~��������u��/��	���Ʒ2�v�ɽ�*<e2G7���7R��ɽ�*<eɽ�*<eɽ�*<e3��$S��x��kNL�0�ۧ��5�a⫏�x�bb����G\��}�}k����4�����l�G�䗴W�����ɽ�*<eɽ�*<e�VJUT���T�$�KU)Bf��S�H}Wf���̃\e񧏟5�����Z�r�_`�m���Q(�>·�ۃRIɽ�*<eɽ�*<eɽ�*<e����a�d!p*�~����_B}��Awo��o�9�HF���,�CVE�OjN�[ߨ�����|цMh���Ai�5��;#tMɽ�*<eР��
K@m��=V�����t��h�����X�hI�
�U�͵�R}����K���3��n5�!������n�����6�Geɽ�*<e����n��r-�[jvsmO)ɠo>fa�������Z|��g1	��S��`&ꬶ�R���3��n5�!������n������QFb�ɽ�*<e����n��ra����������b'!F�+ ��-�[jvsmL���ǅ�\��}�}k�}	�oK��t�e&5�w��=ξ�ֶz�A>υU�%ߏ�VJUT����j\ܤ�"�M�U�帶Ԃt@��@Z���ŗ��J�pJ��AD*2�&I&ꬶ�R���3��n5�!������n��������d<�8��ЎK�����n��r-�[jvsm�����d<�Ju9���b���4���w���x�򠽄��d<�xg��r��*�zN�������Ef��&t�e&5�w��=ξH7Jq
�8��ЎK��VJUT����j\ܤ�"�V��P ��Ju9���b���4���w���x��˃�6��Rbo� ���&ꬶ�Rb���4��r}�<�P�p7R��ɽ�*<eɽ�*<e����n��ra������0�:@	��0�ۧ��5�"W0�Ѵj����z���͵�R}����Kb���4��r}�<�P�p�S�P'qɽ�*<eɽ�*<e����n��ra������0�:@	��O)ɠo>f;�3-�QZ�H[�MF�z�s]eNN`�CVE�OjNh�����nŶ~m߄�7X��q�ɽ�*<eɽ�*<e�ď����1֬��yv�F�W�����[�A���Pt������Awo��o�9�HF���,�CVE�OjNh������3���$5KG5�td'����}g�ɽ�*<eР��
K@m��=�s�VǉzLS��	�!�(I�Ȏ��v�Oe���,�(��Gt�em�B���&��r>��CVE�OjNh������3,e������<���^�� �R��;ɽ�*<eР��
K@m��=�s�V�/�܊���K�am@��e*��i&1(�J��tL:W�xg��r��*�zN������V̴�c䙈e/'��񡹟��n����!f�� �fɽ�*<e�VJUT��ȵ���� �Ys�Mz��0�ۧ��5�3���T���w���x��bb����G\��}�}k��a1:`-e�e/'��񡹟��n�����6�Geɽ�*<e�VJUT��ȵ���� �Ys�Mz��O)ɠo>f��x����Z|��g1	��S��`&ꬶ�R"W0�Ѵj�/�����¯�>�Pp传]�RH�ɽ�*<e����n��r��x�������b'!F�+ ��;�3-�Qm�њy:~�9�[�P&ꬶ�R"W0�Ѵj�/�����8t��4hWV�!�(I켚<dz�Ui����n��r;�3-�Q<�3�N��!�(I�8�>��z�Oa�U�^�\L��f^b�!�(I�o� ���&ꬶ�R"W0�Ѵj�/������_��`���K�am@���h�n�g����n��r;�3-�Q���/*� ��K�am@��%��K���@Z���ŗ ���Ig<g���4�Qp?��y�ճ�袣G<_B�@Z���ŗ�$@�՛��z�iU�}ɽ�*<eɽ�*<e������Pt������91��?���w*���}.��.�J�}��ʶ��^��p�"��Oa�U�^�  񌄮������8�:�ɽ�*<eɽ�*<e��s '�&B����3�`yxvi!\J�)޺�sJp�<fq9�z�s]eNN`�W7P�%Oa�U�^�nŶ~m߄�7X��q�ɽ�*<eɽ�*<e��s '�&B������@&(�v��ya����3�SF�ɝ[:~�9�[�P���K3���T��r}�<�P�p��K�`�W�����ɽ�*<e����n��r��x���0�:@	��,�o��v����M	~c���ġ�H�q/��W7P�%Oa�U�^��3���$5KG5�td'����}g�ɽ�*<e��s '�&B����3�ǉzLS��	�!�(I�8�>��z�E��+)S���!�(I�o� ���&ꬶ�R3���T��r}�<�P�p�"vЅ\�����}g�ɽ�*<e����n��r��x���0�:@	��˃�6��Rb8�>��z���V(���D�K�am@�&��r>��W7P�%-�j�L膲~���˫+&\��p��̵��F��X
ɽ�*<e��s '�&B���i��.�*��w�U.4��odI%C�2g#9+��dK'mgS�}!�Lڜ<��q��M��!Ae��q����C�輒�b���X��j�x"x`һaB�ɽ�*<e[���g�Q�|�������\�����w�U.4��odI%C�2g#9+��dK'mgS��n �u�HYz�s]eNN`�W7P�%-�j�L膲~���˫+���TiIAв�2Gɽ�*<e��_ގ�|�-��(I�z���� ��W��Ľq�>	����I>/�4	��,���/��	���Ʒ2�v�ɽ�*<e-�hm��>0����/B!V'Ba6j�^�T��ɽ�*<erL۪w�Ib�(�틪���]�b�^�!]�?T�R,�&���q�.��W�b���4���u�6����k�~��j�蕘��:2�ξp�޳���~�H����uŬUg/�Qa,�ߴ0�Aw8��a�pN��.��W�3���T���u�6������W��
ē���u��ċ�LY-.fL!�7���U��?Ӊ�xCm�D���X��X����#�Q��/!M_[VǮ���D������q�7᳁�#h���VC扢 1�l�����͏b�^�G�uT��3�&�wU8���-ޝnH]��<�"�".$�B|�G�v3<���@%�BM���!8�r�.X�'~�;.N"��yfs��	`���
��?��!��>	|�W���@F0�b�(�n���8E��T�bP���]�߰5�;�qJ�~<�Pu_^�=�A�y'Xƻ�2������"�lAc�ڵ�?��'����)ؒI
������{���O;�� �m�ۓyP��y��)zr�k&����J?�n=�l�c�I������#/D^PtH)�|/L�$ɠ_M�x�蹹�Hl#[ė���D�h���\�����eO��y� ��W-sD'�4tꦘ���R#l���w�%�<&qj�Iؾ��$s:������8��^R�������߳�_ەU�6����7
�E�Yؽ�&�b!B����Ż�5"rb�R=�5'�x�u)�l����Xp���l��)c��&pW�,��I�\}��Q�p���w�a�yuB��5n<l-�+͘3+1/�s�<���U�P�o�P�[�omK@�Y���V$���`i���8V�����6~8� VQT�!��t̞�����a�}[�t9ƙ�]�?M=�R�i%���XǮ�O��L$��F*�T��'�]J0:���Z��C����?���k&X�L��iԴ�#�i��yn��2����h�-��MJє�Q�α,Ɯ�<�-	�30�5R)U����}�<r��̻7$T����p0�hi��j�h��4�ۋeN�b�v�w��b�	a��J�K� 6e�!/��bs� ��#&2Bna�&�Z��Ov� ���Ҡ�;��NE���w.�KL�k���IT��1�&����hx4�.�2w�C����p~rևb?@m̳�x�t�e-GT�)�q4X,���;�l�@�i"�^�n�؂�#����Xp���l��)c��&pW�,��{i�������K���������4\��]�찴�}0����[P���Q�P��b=��K�X}(�K�r��������gND��7ɽ�*<eB�j�^9�6�v2�gU0)I�P�z\��Ur��D����`���ڭ�b�o1�`oXK��,{���,+�ۘf�hAU6]?�7e���5�_�@[;(�|Ͱ��J�kpa_��Nɽ�*<e�ߐuX�q����h��pɽ�*<e��U�ۄ��2��t�f^�䍣��ɽ�*<e=e��"�5%�!���P��mr�B�j��O\��v��o�z�Z��6�;���ɽ�*<e�
v�ƒm�9(ύ��Bɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R鴼�+��,�����]��ƚ���ɽ�*<e�Xꦻy~�q�����e��1� �����Ŀ�O��h
�K=4,4���?w�,�"�m� ����F�i���!`��Y9�SGiWw�!I�2�١���]����~�H����uŬUg/�Qa,豄T`���/����?�(<����=	5M��%/vZr���m�3'k:�4Wu�?X�g�-�n��qE�����4u�
d��R
�W���d��ٰ#s�V�� ��ɽ�*<eH�*��h�A�B�R$ \�^p�!P$����sb-�j�L膲~���˫+�a������h
�K=4ɽ�*<ex�\�u�p\�Ì�ut�RN!ŀ٣O��Z����P���'�	���^;���^�f��R��IITwN%@QQ�]�Q�Mɽ�*<eNM{9q��ɽ�*<e��_NN�ήG��q���Su���eD�r�U=Y��t�t��ͼBoO��B�Av�'�Bɽ�*<eɽ�*<eҝ[��R�ɽ�*<e���$�*��c�q�΂5�7��dhS*��j��)�o���=��-l	*vɽ�*<eɽ�*<eɽ�*<e�}�F�IH����H���H9��Y9�SGiWwSu���e˴w���{�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���8�9��J��V�B�fd����r��..+`��i=�Z ���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e����<T���Lc ��Z<|Y�M�U�帶�9)�c�d�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e_e��U������ѩ���c�nF�ʔ1�/���%��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r��=�wYh�ǵ�L�Y��6_�DhY��F�(�B)�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���8�9��J��V�B�fP��옸�z�o����{��Q�h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����<T���Lc ���O�	����Ъ�<F	���t�nj�'%萚 tɽ�*<eɽ�*<eɽ�*<eɽ�*<e_e��U�������i�|���}�3|wU���/���%��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r��=�wYh�ǵ�	�P"��49�iv ((�B)�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���8�9��J��V�B�fP��옸��V�\Y�L���{��Q�h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����<T���Lc ���O�	�������$�	���t�nj�'%萚 tɽ�*<eɽ�*<eɽ�*<eɽ�*<e_e��U�������i�|���}�[M������/���%�ȣleg�׿ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r��=�wYh�ǵ�>�Z�('ߛ�M��8�(�B)�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���8�9��J��V�B�fP��옸��a��vQ���#:X�m��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����<T���Lc ���O�	��	b=�(|�4����8�F�'%萚 tɽ�*<eɽ�*<eɽ�*<eɽ�*<e_e��U�������i�|���}��n�[�����At�;Ӷȣleg�׿ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r��=�wYh�ǵ�>�Z�('�}{p�'��c(�B)�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���8�9��J��V�B�fP��옸���vX���#ۑ��th�h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����<T���Lc ���O�	��	b=�(|�4�6;�ɰv�'%萚 tɽ�*<eɽ�*<eɽ�*<eɽ�*<e_e��U�������i�|���}��n�[����-��р�ȣleg�׿ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r��=�wYh�ǵ�>�Z�('�ˍ�����(�B)�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���8�9��J��V�B�fP��옸�I�rJ���͎	�&���h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����<T���Lc ���O�	��	b=�(|�4'X�NJ���'%萚 tɽ�*<eɽ�*<eɽ�*<eɽ�*<e_e��U�������i�|���}��n�[����L��43��ȣleg�׿ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r��=�wYh�ǵ�>�Z�('����D�0��(�B)�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���8�9��J��V�B�fP��옸�꒩V �x`���nx�h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����<T���Lc ���O�	��	b=�(|�4����8����'%萚 tɽ�*<eɽ�*<eɽ�*<eɽ�*<e_e��U�������i�|���}��n�[������܈A<ȣleg�׿ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r��=�wYh�ǵ�(M��䔸�
尌��,i�;��h
�K=4ɽ�*<eɽ�*<eɽ�*<e�VJUT���8�9��J��V�B�fP��옸�G��[��i=�Z ���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e����<T���Lc ���O�	���H�-G�+�e��>� ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e_e��U�������R
�CI���� g�+�����ʠ��6���q|���ݓ`���9n22r�h���Ɯ�h ʋ 2N3J���ɜE.'ѳ��w��ǋ'H)�@wV]��%�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�s�?O��oaf�	��,Jr��v@�0��BkJ&�(�z~�(�^(�~)�����p`�ժH���ɽ�*<eX���Ѯz��<I}�����$�Y��# N��������l�m���t�Yc*��\P�������%�8�v�r��?��&X�o��*C���w9:;\B���١���]����~�H����uŬUg/�Qa,�#z�'�?ḑ��g�DAuUI�,-Я���q���<�����_����Ctb %+��t�s1�Q�]�Q�Mɽ�*<eɽ�*<e�R%�1�Z�G��θ��x�H����Z@�a8���~��91��?��M
����ɽ�*<eɽ�*<eNM{9q���Ef�]���̲�E6�-G��2���3r9$6 &~�!�*�X�����s�ɽ�*<eɽ�*<ex�\�u���U�&4�}p�5ĕr��X��\��g�����6��n��_Lq f�&�������Y���:cl ��C��z󚅔��Q}���5�lcnNMG���뿓�ح׽��J�OK|��Qڨf���xɽ�*<e��Vϣ��c��#�����	/���U�ۄ���d���/)��H/��ɽ�*<ed��Ję���'�D&����A���U�ۄ���!���7�%�&�����V����Fd��Jęf5-�M0,�3��x�K��N9�-(�/��!���7�%$�A��˼����%�G��4��Wzhp�I�ۿww�佦i0Oh�!���7�%1�@ͫ�����e�ʝd��Jęs�Ϭ(�����Z){Q��r��<�-<n���S��̹尮l;�DhY��F�ɽ�*<eg��1-P���h
�K=4ɽ�*<eɽ�*<eɽ�*<e�����^��
:�*�~�sh-�ߠwo�	h�["�Y�n���(�틪��>U� (85�׻\-�!���-l	*v,4���?wL���xr��<I}�ԩ6�ֺ6��b��M&[)�i�����3r9$6 &(d�!�\U�>:�ɽ�*<e,4���?wɽ�*<e�w��ѹ����)��Y�q]�iʳ1s]u۷�ܓ���u���$@�՛�f��Iă�Aɽ�*<e����n��rɽ�*<e��_NN�΢jET�%���:��*�s]u۷�ܓ���u����Q(�>@�ࣨSɽ�*<e����n��rɽ�*<e�0�i�X�wb۳.��:��b��M&���kp��^�� ���y�����ɽ�*<eɽ�*<e����n��r���&B��G��θ��x�H�q]�iʳ1��~l���zG����}��h��ɽ�*<eɽ�*<ex�\�uɽ�*<e�m=����9í�>0\͟�:��*ȟ�~l���G�e�2� ���9�^8�7ɽ�*<eɽ�*<ex�\�uɽ�*<e���$�*�u��|���-Ȳ�N�#sAyA/��6����[ɽ�*<eɽ�*<eɽ�*<ej	�%w\������~�W%8n�B�K*�]�ɽ�*<e(�B)�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eu;�Qݷ�2U���m)�[��mk��畬��+ �0��MK�s�Zɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곑f�[��!<�ɠ)�Fi=�Z ���ɽ�*<eɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ��`���)6�LQ{D���b��M&ݭ�:nB�r/eJR�k�/eJR�k�/eJR�k�ec�*�S�ŧ�s��Q�V�B�f�]&��,�gj�T�1'�� oحɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�����/�\U9��8P�|�� ����!i�#%}ʔʵ�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��M�R��Lc �<gcp2�Š����d<�- �Ƈ���ȣleg�׿ɽ�*<eɽ�*<eɽ�*<e�VJUT���	D��:�^�����%yeTQ}��V8��+ Z���z:�-q26�\�ɽ�*<eɽ�*<eɽ�*<ej	�%w\�����TZm��I����'����V8��+ Z��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<eu;�Qݷ�2U���m��̲�E6�˃�6��RbH�a���akQ�]�Q�Mɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ�f���t��(yaf��ٿ��{��Q�h
�K=4ɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ��|�KLǍ+�����&ɽ�*<e�����l�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�f�S�{��%�u�d}l	���t�nj�'%萚 tɽ�*<eɽ�*<eɽ�*<e����n��r�����/�\U9��8P��/1lG%iP��[P�^1�?q�-ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��M�R��Lc �<gcp2��,�o��v�/���%�ȣleg�׿ɽ�*<eɽ�*<eɽ�*<e�VJUT���	D��:�^�����%��`�l{�J�J=�������\	Mɽ�*<eɽ�*<eɽ�*<eɽ�*<ej	�%w\�����R
�CI���$�$�w�'����ڎX����^*<�]�=׺HGh��Ltג$OJ�7��D���c��#���E6�eQp�8R��������U�ۄ��_�P/4c� 0��%rɽ�*<e�/���%��X��cQ�]�Q�Mɽ�*<eɽ�*<e�VJUT���?�(<��ɽ�*<e^��
:�*�~�sh-�߱�e�[v-%�ؽ->*W-�hm��>0����/B!V'Ba6j�sk��,4���?wɽ�*<e@d����і[.�[����n� Z1�o%���G�c�тQ@ަr�����q�0���BoO��B���K�`�h
�K=4{Or,0��"�������j��T�6��V^�í�>0\͟�:��*��w����	�	�hT�� u�W�g����TiIău�Y�'x�\�uɽ�*<eɽ�*<e�0�i�X�^����y�6����-�Dz#A��G{M��u����s��\�gJ�������f��Iă�A����n��rɽ�*<eɽ�*<e�Ef�]���̲�E6��!I�2/��JZ�+�[ߨ�����|цMh� ����Y��\U�>:�,4���?wɽ�*<eɽ�*<e�JLs������̲�E6������d<�"��È��[ߨ�����|цMh8t��4hWV�!�(I�G�;8�;�/ɽ�*<eɽ�*<eg*D����Vm�B��� Nzw��"vЅ\�J3�W�`>+��6�-�^"����Hv���"���<���^#z�͌�?�(<��ɽ�*<e����Ħ�
V8��+ Z�zh#��d��-QJ����&�H�@�p1W:�=����ɽ�*<eɽ�*<e,4���?wc'w�>�~���˫+���"ˡ��LG��..+`���/���%�2G7����ᦲc�ɽ�*<eɽ�*<e�VJUT���?�(<��ɽ�*<eH�*��h�A�5B�	��Y��# N��ɽ�*<e����wEF���R��0ɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e����������BZθs�X��\��g�����6���q�0��?��`����9�z�Y�����Ɯ�h�[�Z�~�q>R}9�܆�h�q+�yp�Dm��j"�Vj�	K�ؕ�U�@>�����Z�'[P�u�ɽ�*<e1? ��6�2��p�ɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e^��
:�*�~�sh-�߱�e�[v-%��1�>,�(�틪��>U� (85�׻\-�!���-l	*v����옙�;��R�˴qZ5�+�/I��/�F�W����ɽ�*<e�'3�FJ�c5U�2#3�^�&��Q�]�Q�M!����M�b�%��)�BoO��B����$�*�%�ܧ�	\�j�<�U�qD�r�U=Y��u�[��91��?��M
����,4���?wɽ�*<eɽ�*<e�Ef�]�ԩ6�ֺ6��b��M&�DD��,�J����3������l�V�\U�>:�ɽ�*<e�����ɽ�*<e���P��Z|[s%�o,�o��v$����sbOa�U�^�(S	�f�w�_jk�#��ɽ�*<eҝ[��R�ɽ�*<e�2R&�N5݄p��P2��࣏�>�m�B����Z�`�n�[}ͣ��T���'����V8��+ Z�7F'�]hɽ�*<eɽ�*<eB��gJ��A���4�Qp?��&�E@s��K�am@��z/����`�@Z���ŗ�Z�9�V8��+ Z�����?�(<��ɽ�*<eP�ay��b���4�Qp?�U�ݣ��d��-QJ��'�	���^;���^�f��R���R�S��� ��ZXd�"�ǳ���r�~���˫+���"ˡ�6�v��������P�$����sb-�j�L膲~���˫+&\��p���M
����ҝ[��R�ɽ�*<e�`���{�"M��
f��S�Hɽ�*<ePer�"��۞�XZ�v� ����Y�^W���}/2Y[v�_�ɽ�*<e+�n�/�G���!�f��=#c?�V�Y���n5�!���S#+�Z��2p[�������Ɯ�h�[�Z�~�q�q��N�S�U��h��OK|��Qڨ������6��x�B��?;�{�,��-soۘ���;k�7�_��g='ѳ��w��ɽ�*<eǋ'H)�@wV]��%�ɽ�*<eɽ�*<eɽ�*<eNM{9q��:j���+�oaf�	��,Jr��v@�00��� �<���^�jT(�z~�(�^(�~)�����p`�ժH���NM{9q��L���xr��<I}�D��݇�3�W�D6�fɽ�*<e��ۦx�/�����¯�>�Pp��9�^8�7,4���?w��!�2X���d�'\�����Ş��i91��?��Nd"�O���xM�Aw�i�e/'��񡹟��n����AE
!�ɽ�*<e�����ɽ�*<e�m=����9o;���5���������ƎAXU߮�MLŞʅ]]�����>�Aft3�ɽ�*<eNM{9q��ɽ�*<e�� Qx�����,}�k�G5�td'�{�������&k���˱M���ݾ��*���F�V8��+ Z�iE����nɽ�*<eg*D����Vm�B��� Nzw��"vЅ\�J3�W�`>+;�3-�Q������I7Is[���V8��+ Z�7F'�]hɽ�*<e��#)ϫ��K�am@���V���/�Su���e�/���%�a�������'������W:�=����ɽ�*<e����n��r��݌�</<_�BU	���v��J�};\B��ɽ�*<e�sĸ(�A��c5U�2#XEߵW�,Q�]�Q�M�VJUT���?�(<��+�n�/�G���q�����`�2�ɽ�*<e�z?,�y��u�[����l�G���h
�K=4ɽ�*<eҝ[��R�ɽ�*<e:��8*$7�K�K����̸B���=RMq��-��@Z���ŗ j��c�̸B�����y���C�NM{9q��ɽ�*<e8�q�ѱ�V8��+ Z��Moi��v���<���^"*��g)x�h������3,e������<���^��y���C�x�\�uɽ�*<e����Ħ�
V8��+ Z�"#��K�d(T�F(��@�j/�j���̩;IJ�}�o���ɽ�*<eɽ�*<e���  I·�#=�Ԣ�¼�(�!� 4���:o/���?��ɽ�*<eS*��j�Ǐl���SI�\U�>:�ɽ�*<eɽ�*<e�����ɽ�*<eD���p �W|��C���Nd"�O���/���%�.�6�o�&TD�>蔽iɽ�*<eɽ�*<e����n��rɽ�*<e!�T9�u����Nk�QWk�HZ�ɽ�*<e�������k;c���xɽ�*<eɽ�*<e,4���?wɽ�*<e��vVK�`���;�	Ei���!�)�49�iv (S*��j���LQ{D��y�����ɽ�*<eɽ�*<e�����ɽ�*<e�4ł���:��������9���wo�	h�[��������rq��&�������ɽ�*<e,4���?wɽ�*<e��vVK�`M�L>�;>c�'�i���臰z�IYLy�q]�iʳ1�������/���?���AE
!�ɽ�*<e,4���?wɽ�*<e�H��g澁_d�Ǹ��#��6*+�'���g�#w�'�S 5l�S*��j�ǌ����6�%��;�	bɽ�*<eɽ�*<e�����ɽ�*<eVd�����	�3��c� g�+�����ʠ��6���q|���a������{�� ��5�ג$OJ�7᳋��(�4��mq2����Z�'[P�u�ɽ�*<ew�;L�::^�Q��	�ɽ�*<eɽ�*<eɽ�*<e,4���?w�4����k���A�X:蝖`�uɽ�*<e�Xꦻy~�q�����e��1� �����Ŀ�O��h
�K=4�}�F�IH��, ��T�ԩ6�ֺ6��b��M&/��JZ�+�[ߨ�����|цMh� ����Y��\U�>:�,4���?w�&X�o��*C���w9:;\B��ɽ�*<eQ@ަr�����q�0���BoO��B��ᦲc�ɽ�*<eҝ[��R���_NN�΢jET�%���:��*�Dz#A��G{M��u����s��\�g�l$aw"@�ࣨS����n��r!�T9��v��J�}���:��e
ٰ���˫�Q@ަr�����q�0���BoO��B�"�#F��8����T�ҝ[��R�B��gJ��A���4�Qp?��&�E@s��K�am@�{	:ܢ��l{M��u����s��\�gI7Is[���V8��+ Z�7F'�]h��#)ϫ��K�am@���V���/�,�o��v�/���%󬭠6�-�^"����Ŀ�;3:-��_jk�#���VJUT���uUI�,-Я�ƚ��wb۳.��:��b��M&Dz#A��Gm��=�s�V�����l�V�\U�>:�ɽ�*<e����n��r\/l�<�]��<}�l=2���mɽ�*<eA\x/~�!r}�<�P�p�ᦲc�ɽ�*<eɽ�*<e����였m=����9í�>0\͟�:��*��w����	��@Z���ŗ��Q(�>@�ࣨSɽ�*<ex�\�u���U�&4�h^�!�����ym��Aٰ���˫�A\x/~�!r}�<�P�p"�#F��8����T�ɽ�*<e���������o���S�B���@%;�� ����K�am@�b���k�k�@Z���ŗ�Z�9�V8��+ ZL�q�e���x�\�u����Ħ�
V8��+ Z+�+o��[}[��z��I-듈�<���jA�ԁ�@Z���ŗb��i���sX!���x���+�v�ƶ2�]�H۝�ɽ�*<e�
v�ƒm�9(ύ��Bɽ�*<eɽ�*<eɽ�*<e��:R�XE�&I��}�, ��T�ɽ�*<e8u�U�'\X�aҥ��|2R+%�~�!�*�X�I�� �p�Z���-\dE,>������D\ȯ��!I�2�/���%�;�3-�Q������X��j�x"�&ZReX�����n��r!��2����jN�̓������P�ɽ�*<e��ۦx�/��������Ai��h��,4���?wW���P�#��6*+�'�F�W����ɽ�*<e�xM�Aw�i�e/'��񡹟��n���W:�=����ɽ�*<e����옫��$�*K�K����̸B����eK�ֆMLŞʅ]]�����Z�ͥ�!yϦM�|.,K�%-
+[8�q�ѱ�V8��+ Z��Moi��v���<���^��5�����,�v��l�����z�n�yϦM�|.9�<7�������Ħ�
V8��+ Z��̲�E6��!I�2$����sbOa�U�^�  񌄮���y�����ɽ�*<ex�\�uD��N_��^[V�Cg�����P��/���%���x����'�������AE
!�ɽ�*<e����n��r�`���{�"M��
��U�����ɽ�*<e�'3�FJ�c5U�2#3�^�&��Q�]�Q�M�VJUT���uUI�,-Я��`K�f��9üI`�̸B���w}TڽԱ���u�[��{M�y0��bm�B���m�����ҝ[��R�B��gJ��A���4�Qp?��^� |����<���^KK1�3�����3����^����K�am@��m�����Y[v�_�P�ay��b���4�Qp?��������Jd�q/��DD��,�J����3����\�
p)�1���ɽ�*<eY[v�_�
�'63���������$�$�w�'� �۟�6 �D�G�9#|�����N���Q�)y��$�-�bJ	��$�1�x0Ycɽ�*<e�%�G��<��;τ��2������7a~�	��1�z�'G�7�߰XnVC4[!7,���f���xɽ�*<e�:�<�.�ؗ���v��_P!_��~��7�q�Xm.��ߐuX�q�g']5��kLDQǺ��@y~�^+���B�j�^9/-E��+lJ@Ҷ#�hMU)�_>%"	�E׋������z�{Ά�[����;(�Y�>���?�L��P�a��D��VZF��m���|(~��
��ߐuX�q�����V��U?��4���[���A�.���)V�T(�<7���_P!_h�Ү����U��h���Lw��g']5��kL���RI?��U���v�L��P�a��D��VZF��m��-��y�����ߐuX�q�����V��U?��4�J�����.���)V�T(�<7���_P!_�6�̚r��U��h���Lw��g']5��kL���RI?��g�.@L��P�a��D��VZF��m���LD��@�ߐuX�q�����V��U?��4�H���.��.���)V�T(�<7���_P!_��6��kP��U��h���Lw��g']5��kL���RI?�����X0�L��P�a��D��VZF��m��V�D�����ߐuX�q�����V��U?��4�sXi��L�F�.���)V�T(�<7���_P!_̅�k=�g�U��h���Lw��g']5��kL���RI?�)nV�i�(�fkN�F��&B�B_E�U?��4�*��@M�aU{� P����(�틪���fڸuO��y'p�k�&��중���{}�gn(`m�R��y���C�ɽ�*<erL۪w�Ib�D�4�i�K{��%B{$'ѳ��w��ɽ�*<e��=!��(]��s�kɽ�*<eɽ�*<eY[v�_���ܑ��h"z<�'~�V'Ba6j�"�Y�n���(�틪��>U� (85�׻\-�!���-l	*v�}�F�IH�u�c�W<� ������,��V�X�˄����pɽ�*<eɽ�*<eɽ�*<e�VJUT���	D��:�^�����%Jr��v@�0{��Oũ�&(�B)�ɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ���m��&��7�H.�M	���t�nj�'%萚 tɽ�*<eɽ�*<e�VJUT���	D��:�^�����%Jr��v@�0z�aN±�(�B)�ɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ���m��&�~�C(	���t�nj�'%萚 tɽ�*<eɽ�*<e�VJUT���	D��:�^�����%Jr��v@�0%�ØX�h'(�B)�ɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ���m��&��Ҧ�d	���t�nj�'%萚 tɽ�*<eɽ�*<e�VJUT���	D��:�^�����%Jr��v@�00ƶ��le(�B)�ɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ���m��&��B:�F�d	���t�nj�'%萚 tɽ�*<eɽ�*<e�VJUT���	D��:�^�����%Jr��v@�0D,�.�e(�B)�ɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ���m��&�}�Z,��g�	���t�nj�'%萚 tɽ�*<eɽ�*<e�VJUT���	D��:�^�����%Jr��v@�0��ܕ�=}(�B)�ɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ���m��&�{(��V��	���t�nj�'%萚 tɽ�*<eɽ�*<e�VJUT���	D��:�^�����%Jr��v@�0+"��B;(�B)�ɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ���m��&��w< �:	���t�nj�'%萚 tɽ�*<eɽ�*<e�VJUT���	D��:�^�����%Jr��v@�0�F��=(�B)�ɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ���m��&���Z�`��	���t�nj�'%萚 tɽ�*<eɽ�*<e�VJUT���	D��:�^�����%Jr��v@�0�x�6Kx�(�B)�ɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ���m��&�9f<vR� �	���t�nj�'%萚 tɽ�*<eɽ�*<e�VJUT���	D��:�^�����%Jr��v@�0����8�(�B)�ɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ���m��&������*	���t�nj�'%萚 tɽ�*<eɽ�*<e�VJUT���	D��:�^�����%Jr��v@�0�0
�d\,w(�B)�ɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ���m��&�8K:5���	���t�nj�'%萚 tɽ�*<eɽ�*<e�VJUT���	D��:�^�����%Jr��v@�0��Z�1��(�B)�ɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ���m��&���*�r�_	���t�nj�'%萚 tɽ�*<eɽ�*<e�VJUT���	D��:�^�����%Jr��v@�0��b�Ǜ�(�B)�ɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ���m��&�i^#w�)	���t�nj�'%萚 tɽ�*<eɽ�*<e�VJUT���	D��:�^�����%Jr��v@�0٩���Ò(�B)�ɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ���m��&�Ѣ�yO�	���t�nj�'%萚 tɽ�*<eɽ�*<e�VJUT���	D��:�^�����%Jr��v@�0�
n�z49J(�B)�ɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ���m��&��Do.��	���t�nj�'%萚 tɽ�*<eɽ�*<e�VJUT���	D��:�^�����%Jr��v@�0.�^�<�eUXec��
ɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ����Ve:}Rk!��^�(
P�����Wm��:Y�f�H3UU���f�O@g�IFS�w�s@�����4�
�����%nġCB�I�t�`H�Q����U�xl�(T�W#�(�*� �.6p@�*3d�#_�0!s�,�	���
6�.8�0�T��(�H���-)�|�d!d�H�d�h�ݔ�x��{��õv�̟��������.s����g ��$�L��ow(7ALۗ)��/��	`�)�h��{̠����Lʉ/[¶���`���c��� �	[�w:���ע��������t��E�̎����D�<L}ڈ�����dn'y&���3��ͨL���K��a9q;���]��e�G<���ߤ#����ө�((|�w��M{� C<�ls���|����䋇�æ��tg������a��4W}����Y[A`�_Z_MyV<tn�||oKװE��"
8��o���l��͡U�R�4�t���#,�>�Y����,�:�+[��epՈI��	n��WO�.�<8��]���f8��H�\J����K=҉7�#������g~�nR�&x��l���Hwa_i��\{��ЍM�Cʌ���H�v���5������A��\��G������Oc]����s��� �F��.�8X��)8�\/,AܥЍ�ө�	I�\���YVeX���V�E{�49��������4�=z��F		DAu��6YhzoC-x�i���
V�r&A�V�6�.j���|R��Ǥ_�|�P��L���Xj��)�*��e/6�5��0�u�rq���	�//:��;�$S�,9�{M���S�w�s@�����4�
�����%nġCB�I�t�`H����N�,9�{M���)_d<�cYb�'����4�È}����Hc�;�Y^�U=���8��u������Qk4]��
�k���_=������Y�"�WZ9���u\�a݀P�!s�,�	���Π��U��~Hfu��Ԯ�΍T�:��S� k/!M_[V�I'�
n� 70^�d�e»�-0^��,�:�	S�uP�M�zK!�g٪�'�)��F�p�	_ى�#�9�$�oWU� ����L�m�C��#��;����B�	?�gwC�N�O�lK���K)��F��P������_#Ǚ��R�����'c.�	?0-� ����Jv�T�`���LZu��,�K���G.|DT����(PЎ��=H��|�j�U�d����q��0S�tO��t��t%~���L��b��+[��epՈI��	n��WO�.�<8��]���f8��H�\J����K=҉7�#������g~�nR�&x��l���Hwa_i��\{��ЍM�Cʌ���H�v���5������A��\��G������Oc]����s��� �F��.�8X��)8�\/,Aܥ�1@U�����7�Y�}ފ	�=��ϝ�p:�A �Ы���VI#�1z���x�q��Ǝ�b\[��½�#��$̆���5��0^v�'-�r�D��6�^i~��b!�t�&��9W������U��!��?�0.܍�G.I�TVzin:+�w?�>�X�L�7����=pS��-�qS�*':���-,;m_��Dȫ+@-p�\kgd\/��~�d��yA�/I��d�H1�J�K
5�������iSUk=�Pq�vGfG�/1�l�[#�e�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S�`�	�hY�*L�2x*���L"M��Qp�wW��-4০F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��"�iS{�؛��}snv2��z��b=�D2�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S�X<��a5���I uA�6[����S�2͙gG�7W��d(�e��'_>g�Q]e8�3�F�ڄqÖ��T�̡���C�O	����]�ͻlU��5_�rG���-��V  �쵶6�1?*�k+�*FƠ�h��^1_�}J׃���2�$D���Wѵ/5�gD��mv�Bӝ`Y7�:f��$Cl#�8H�r|�C��� �y��ug�s��^Jx�66:��b� z5��ɽ�*<e�ʻ�;)n�wa�.�g�ӳ�q�s��^Jx��h\��"r{��Bd�ɽ�*<e���=s� HK����6�͟^ɽ�*<eX1��rぱ@��Z�ݐ;��?t���C��4�L�)� UPWd�}�q�80�L^ʔ��Ɨ�̜�X�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8���j�o;��ph9!�4�hԚԾ3�81R�c���E�zַ���@B1Y-�q f�&�.�����j�B;ߐ��yם�A�<�Ʃ6��/W�����a3m����@����xw��E.8Ԙy�9ɽ�*<eƚ������=��c��v\�I;����u8�X�J�X���	�t�k�(IZ��ºS����3L,Ch�b> |�!N��� ��#*ɽ�*<e��݌�</<G5�td'�fwJ�W��5����_k`ɽ�*<e�*�S� V8��+ Z ��ϫ)��;��t�^	�'E���.�^<�
:�ɽ�*<e�C�.��Dt?�Ѳ����9��ɽ�*<e[����Eh{3���
����9�֭�OF���c]ǻ8_!���kJ��f�[>���ɽ�*<e�g?k�Vtև̸B���95tH��f�[>���ɽ�*<ee&����h�V8��+ Z�40�U�a���D9$�UQ�ʲ5����_k`ɽ�*<e>"��;a��I��&6=��^���Gg}4���R/�B�a�h�ɽ�*<e|"y�׫&��r�� �%�]'E���i)�7h���Ɨ���#�����F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�ol&���rl�8ko#'DV�X�^�˪l�VUQ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q�݂���q�EĄ�#���&�|�D�µ��g���>��g]�?���'{�5r{[����Eh� ��̭.��>��������&B����!2��Ȝ��X|�YA�Y��g{M�y0��bm�B����*�b���G5�td'-�f��ݬ��!�2X��˃�6��Rb�����E�"vЅ\�"�1K�;��]�P�.�F��K�`ƞ�rL�mD%��9)�L� \f.��_�rҦ�S"Rjm�@^B}�/�x`B�*���8w�PO��Y���X��k����˾���=O��E�¬뤴��RL�-s��2[��xZ�ݑf�v�t-ձ�b�9�5�ҹ��m�]�!�m,�H��B".��K�`����K�k���,(n]�P�.�F&��N�����8�!�|����n��r�w;$�y�%��$>��v�I�pKP�7ٝGy��v��,��}Rk!�:�ѾM ~��Í�a�h��?�9���ْ;0b5��u|R�2�i1���u�\��u�t���JX�o�'���tM#�/��t'���hX�O@g�IF)_d<�cYb�'����4�È}����Hc�;�Y^�U=���8��u������Qk4]��
�k���_=������Y�"�WZ9���u\�a݀P�!s�,�	���Π��U��~Hfu��Ԯ�΍T�:��S� k�7��`x\ `L����JmB6q~q�~�i7 :���Iy�;�nų�j �@V��"WP{Y�GT���8�Y��i����QQ*rbH�iA�UAKTnО�>����x�})I)���()�6��9w嚋.�����_xUʯfK���� �]Ե�:i��Ly�|y�ި���6�ʈ����I_�Ut�)��7�џ�q�s�Mv�'��X�)����qӬ�\ԗ������nx�I��	n���#���o�oi�8�,����̜�ߑk���g���>�0 ;��od<~R��Ǥ����e�9�\?%&�/�~=rN��uL�7d̈w�U���YEL8��L�Y���ay\�n ���J?|��'�[����K���3��h�A5�oD����S�_>gN0e�,F��Т�����[���ɛJ�z6Ǡ�&�ǅ���7�Y�}ފ	�c����$���D����,���AI'�Q�Oﴽ���������
����-��
�=��U&ʀeH��J�	�5!�`G$j`{�+!�Nh�z�{&�@�E�� �/.�:Y�f�H��� �� �&���2�i1���u�\��u�t���JX�o�'���tM#�/���g���x �&�����GX��a��Xڟ3�8�H�d�h���� I���}�t�wI'[]
*�J���oE����:��C�$k5p!,�7ڐ9� ��h��'i沃�Z}����Hc�9�%�\T|Aů� �B�#��t�(a�������bc+Ji �8s����6e���%���2"��
��4N;L�Oc]����m���x�?���wIF��E��OU���2ޔ��e�����{�n�q�r/<��\�D?('h(�m�W�K.j\�NIf���'Q+j���p�D;&��'��K�����c�׈�}���	'��@Ybs����Q��� ��ɬw��2,mD9���\��w�0��8w���c�Y�l�%�tB�;��Ha�L�zַ��-ro��S�7>�<S@��9jj ����̜�ߑk���g���>�0 ;��od<~R��Ǥ����e�9�\?%&�/�~=rN��uL�7d̈w�U���YEL8��L�Y���ay\�n ���J?|��'�[����K���3��h�A5�oD����S�_>gN0e�,F��Т�����[���ɛJ�z6Ǡ$^�H�#��]G� ��\J���H�����v\�k�tf�����0U������J�yP��}H�{_�.�@)1�7-��H�&��_�6�*�q#�L
2�������̹�"�j��;�kԐH`�Q�����p��N����:��*D�)�=�����ٿ+��Cs77v�������%�mv�Bӝ``�PF�B|O��$����tk���}Ո�,�AQ]�h�j�v���� ��=?C�eU�(p�a�܂�&�>\���;�;���L�H�ZoF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�8�v�_�m2��h���9'e���)�nTz�144zO���=X�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�4)�}Uh���"ﾆ��ъ��>?C������F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�$��0ƺ�R�f
���Y�p~rևH���Nv��7�:��E�fV�,��G�VF�Ar��hԚԾ3�81R�c���ۆ�28� �@B1Y-�q f�&�,/�z/�sw����P�K��3,�g�ӳ�q��.�"3$��&&�����m,�̿ŕ��C4+n��ʌ?a���W�-b(g���⾟�i�,z��x);���o_���W�[�Pp���&|R����h$@�E���wɽ�*<eJ�N�B�%����GO��g���⾟��/s!_ǁ;���	���V=�"�ɽ�*<e��g�E����h\��"��##<�Zɽ�*<e���=s�e���82����ӟ�0�ɽ�*<e�dcL�+C
(_?���#��b��s�um$E��hi�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8��O>3���UW��]T'3���^��w`؟Lk�S,P 09���u�[��b=��K�XG*0=.��Y{79���;��t�^	�SY�A8�f�[>���ɽ�*<e�F�W�����Q����Yɽ�*<e�&�|�D� ���	/��� ��#*�ƞ�ʻ�ܻ�r�i:Mk�F�j4�.�^<�
:�ɽ�*<eXV_�v$m�B���`~X�G�wo�	h�[����@��J��tL:W�s��7ZI��&6=��cf44H���.��|ɽ�*<e\Jԙ�% ���U���������b���>���6��\Jԙ�% �>|
ϒ��ޱ���b���4M�������"�8�U� �n�4�d�FQ�o���������v���ѫe�M�U�帶@3Ƞ�O�����a3mɽ�*<e{M�y0��bm�B���Q�q^P6����a3mɽ�*<etseQ,���F���mI7�;��t�^	�?m�.�^<�
:�ɽ�*<e���!��Uj+���蜵���C��g����{�wo�	h�[vS+ё@|���Hwȭ����O��NH���9c���ġ�e�伸�M*�D��|F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�&���y�����Q��+4�3%�J_�5h�0X�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)X'4M���/v`S^!������F�W���ʲ-�#Y�Rk�\DԷ��J��!�2X��f�2N�2���M`.�A�Y��g��l�G�䗾��ޠ��7�V�)i�g��!^v�!�(I켆����E"�#F��8O�^p=����&B���V��P ��2�>��1���q�ޤO�^p=����{1�o%��w��^��3����&B��M�U�帶�<�+q�@J�F+�m9K0.d�չ�Rhp��Ԁ�F�Y���~N�Ɂ�6�r��s(�?A�Ҏ&�Ё?m�-�,�X�Ÿ�f�2_B@�~%.DI���:��t�%2�/	J��hא�܇*9�2�\c�5��u|R���GX��a��Xڟ3�8�H�d�h���� I���}�t�wI'[]
*�J���oE����:��C�$k5p!,�7ڐ9� ��h��'i沃�Z}����Hc�9�%�\T|Aů� �B�#��t�(a�����z}�E!Ͽ���!Lؒ&�bL�.��. ����lB��,zyj���0_��A�\��B�N��%졖*��j)?��(a�����@��$�G#�ӵI�0��#Ҟ�s�-I@>������BP�\_�0'���I"ʈ�W�rB�������i0aXK��2��H����D���i�6 ��Z�)a��\ `L���c��}W�R�#C,��n�Yx���|��/_��P��r�k���g��� H]K�s��K���{T��
�7`�	�6�#'	��m�:��eH��J�	��[W�DC�"�N�?�ot�'��#~D��\��KB����VL��'�s���7K�f*���b�0qK�s��D�1d�	!4wI�o P��z9����D�����e�mu���H��H�
:��p��؋9i�^��,1DԾ����\J���H�.'a:�s�c�A �Ы���VI#�1z���x�q��Ǝ�b\[��½�#��$̆���5��0^v�'-�r�D��6�^i~��b!�t�&��9W����z��\(u���?�9�o<̀�t����{����f�2_B@�~%.DI���:��t�%2�/	J��hא�܇r���+9}�t����{����f�2_B@:P��dS	nT��e�&��F]�J�������	U�֝�%��LP�b�I�hS\'��/���`b]P�L��ϰ�9_��]-͍)�,\���� I���X�%���=��dn'y&̢���N���ꗳ�)�7��y���#H����^'�2����:W�0s�����S�_>gN�-�:'��$+���G(����^Le�0�[��z����jcbb_�B�,��y8f���B6Km���'�5uEq_�<|7.���|N;X�^�I�[\o|�o�����|"ÝW}�utiO����+�%�Q)=d���E@�׺�F�b3��5����4�fgHg)%�RPz
2����$_�>U�V-'�I��.3	
.5�4w���
ק5�C>��M ˶�{T��
�7`�	�6�#'	��m�:��eH��J�	��[W�DC�"�N�?�ot�'��#~D��\��KB����VL��'�s���7K�f*���b�0qK�s��D�1d�	!4wI�o P��z9����D�����e�mu���H��H�
:��p��؋9i��������a:�#�f"�6]v��P��w�	|"�@Ҍp���O��"P)�6�m�`�� P����Y6Z����*y����,��/�&�5K}�*���ՙ��e'�������s�SŠ��z��Qd_No��H�?&�� 8����y��Z��Vo儢�,)�$����@�H�Z�|�e���&�E�?��`�PF�B|O��$����tk���}Ո�,�AQ]�h�j�v���� ��=?C�eU�(�<�2����&�>\���;�;���L$�����=����H��ºi�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��k^I ��P�u��iXj��a�0�LT�ѿ��3��17�i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8���ա8&�o�	rr��<���b��Pvlu��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�$��0ƺ�R�f
���Y�p~rևH���Nv��7�:��E�fV�,��'_>g�Q]e8�3�F�ڄqÖ��T��N�k|��^�Fϗd��8B`}��z��(V�J�ٛ�c�zr{��Bd˦p3:O�r��E��9��*���s~r{��Bd�� (9��Ơ�h��G7��h��t���g�E��5�gD���9�Y��U�PcY�A X1��rぱŮ�8�5x�*o������,��_dIc�������d�9>؁)#�zNs��^JxMΒ�ӻ�"ْβɽ�*<eN���F<w���P]80�L^ʔ�8ՕmR�%"��jMEf7s�=��4��/s!_ǁ4�W��$��K����������8�Cl#�8H�r�F�W���ʷ��nj;T�E��n�����3�jh��>.��]�u&�D�<��Ơ�h�� ����b� z5��J�N�B�%@.F�rqDZ��F��������sW@k�z$�DS ���i7�%�۞>�8�ꜟ�A�r�J��9W� ��צ^�͌i?���x���,иQ+?�?�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S���S��be�����oz)���ʠ��6���q|���ݓ`���9n22r�h���Ɯ�h�<�ʌ/5����_k`ɽ�*<e�S���H��֭.�^<�
:�����$]�Y�y�Na	-�������a���D9$TRȉ�<5����_k`ɽ�*<e��3�jh���L@(:&��72L%hQQ��p��u��d��)����ޘf�n6�72L%hQQ�E�Ћ��.:����5((яlUj+����1�2P'L�E.8Ԙy�9ɽ�*<e���r�< ��ϫ)��;��t�^	�#�x0U�o\�I;���ɽ�*<e`ύ���#��̿u���E"��R:n0��?�i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S����>��ɝ:������ti<8=�yQaX�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)X��^��6ՊΏ�{��P���c���W�3�cl5�*N�s���M|~�@.F�rqD74������~���P�$�z�s:��7X��q��v����ɽ�*<e��q�Ӭf<ꥴ d�����6�cW�n2L�CA�A~�f���fzP�u��A��'_ؾ�=� j�Z��JПE�[5����[�:��P�~�֡ݻ!�D���8c�@�?��Y�ա|�W2�j"g���fr2�'��2�:@�R���KE�Y�޶���\4�Eۢ�"{�ղ����nUK?-˔ Q�,�n]�"c��\$�� ����%�0.d�չ�R��Q�3����BrW��mVW��c�=O��4f��l�VUQ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q�ݠk��oOLe�fUͪ��{p%WOi�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S�j`▘9��e�=�@侮/�žC
�nd_p�0��2����_��
�cE�H�@~�����"[���0��x�1��2���
�9����C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�HE��޻'�����.в�0q����O ��;���l�VUQ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q��(���|�b��^�i��jP�ab�+�,�!�@�h5m��T�2+��@]�P�.�F&��N���x[���K&��`�7.\�,��2�0���X����� ���/�@���� d!p*�~���iֱ�/5��8��ٞ�bw�x��D��k�N���?���U��r<���QE����r�����׀t���8ο�K����dmk�ג$OJ�7��h�p�4˅��XU�U��q@�+������|;m��v|�YL�ڂ���(|��ڡ��K���"6݋�3���a4�M�Q���X��x�'k��<�D��1�I�>��a��w�����Cſ�y�	�J�n���M������P:խrQV*��\u�Q�o�����q�<��g:�Bح%�R��2Dp�ݏ~�e�ph9!�4�hԚԾ3��Q���d�O��]����;�a��]�ͻlU��Ҏ�_��yMuC�l�g����Z�K�{��ex��D���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<eɽ�*<eɽ�*<e�K�{��e�MO�~I�����1VRKD�vQF��N&d�U�7,?-�Y�������bC�x���b��6�-4�)�_π]Z�$}��b�J�۞F�W���[�&�E�?9D�uǎqh��˴qZ5���JNRy�I�D�J�ɽ�*<e��7�1��W���[�&�E�?9D�uǎqh��gn(`m�R6��P�7kZQ�1	�|�`χ�a$����^�M�"�ds��]W����H9�� �ϵ%[��6ҷ�׸�3�q�w��ΗCf�|����
���2Q�]�Q�Mɽ�*<eɽ�*<eҝ[��R�ɽ�*<eɽ�*<e��N&d�U��j��Eh��!�����y�äB<��{T�_0���ɽ�*<e\���ֻ'���x����9���;�A�-ɽ�*<e,4���?wɽ�*<eɽ�*<eɽ�*<eɽ�*<e+�n�/�G��rq��&�:+�[��sʶ��6L{.���ς���J��^��k)ɬ׼W��#T����i�F�Lɽ�*<e�VJUT���?�(<��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eVd�����$]�7���sʶ��6L&ꬶ�R���J��.�6�o�&}n���%fɽ�*<eɽ�*<e�VJUT���?�(<��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eM��u�^8:���Җ LF�6ҷ�׸�3�q�w��ΗCf�|���P�6;7}o:����v�ɽ�*<eɽ�*<eҝ[��R�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����^��mߠ�]�:.H.�4&ꬶ�R���J��.�6�o�&�_d�Ǹ���ΒQ���ɽ�*<e�VJUT���?�(<��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eD���p �W"!��ٜ;MuC�l�g����Z>[��H����G:fGv�B��-�>�5ɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��r�ό �����B�VT�́s�ڢ>��ڭWH��;��)����&��g��sɽ�*<eɽ�*<e����n��rɽ�*<eɽ�*<eɽ�*<eɽ�*<e��vVK�`^|��]`��V�mB��W�����D}���+H8�|q{+冰�@��M��^��l�ɽ�*<eɽ�*<ex�\�uɽ�*<eɽ�*<eɽ�*<e�@����L_��q���;�d �� �ϵ%[��6ҷ�׸aV�CF�[@�ͽ�Te]��1�k�ɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����^��mߠ�]�:.H.�4��vA�my��Z0B���k�UhU�GG�/���ɽ�*<eɽ�*<e�VJUT���?�(<��ɽ�*<eɽ�*<e1稆���%�I�\�m�ʄ�%�>v;�e�`䷟����{v���)`���#��	�d��hM'��INzW-;�+j8ɽ�*<eɽ�*<ex�\�uɽ�*<eɽ�*<eɽ�*<eɽ�*<e!�T9�u�P�+H�"�o�6�ꪕN#�[K�C:K��.�u�ڇ��C��_	�6��ɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<eɽ�*<eɽ�*<e;K�Raz��|t��{~�y�sʶ��6LTy_2~��	��Z0B���ö���H3�=�Xɽ�*<eɽ�*<e�VJUT���?�(<��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eD���p �W(�$ɯ*���S���)����~�U��ϝO�}�/���>;�# m	�ɽ�*<eɽ�*<e����n��rɽ�*<eɽ�*<eɽ�*<exP�Z�W揔�'��)��] �, MuC�l�g�j7�po�W|9��\�������/���?��Q�]�Q�Mɽ�*<eɽ�*<eNM{9q��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��]/߷�WW���;��X z_.?�P��i�����@�������%�R*
���7ɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<eɽ�*<eЖ��ٿE;i���`C>���z�례݊B�VT�́�Y7W��*�(�2Y�ǫ��8���8��8ɽ�*<eɽ�*<e����n��rɽ�*<eɽ�*<eɽ�*<eɽ�*<e�H��g澚c����2��E+��I�A�hX@��I�b�H汁�
���2Q�]�Q�Mɽ�*<eɽ�*<eY[v�_�ɽ�*<eɽ�*<eɽ�*<e��Z0B��Q��K=Y��I|��w�)3���ӴW��j�1���,�{�����w�9��q�&ɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<e7[��İ���G��͌b{T�_0��ݕ�^6�D���?��B����%O��:��� ���ɽ�*<eɽ�*<e,4���?wɽ�*<eɽ�*<eɽ�*<e�2��9�|�s��
�Δm��ڛ����1V�A`��Cr�W�B�	E�7;	��7�8��P�6;7}o:����v�ɽ�*<eɽ�*<eY[v�_�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e���U�&4�K����!���Җ LF,ҌyX�'�<��|�C�6�vm�y���:��`ɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<eɽ�*<e�W7P�%df!п�jG�7�7�Uz� �[��I�D�J�;�e(<�KB�x�#αh��w$o����� Fx�ɽ�*<eɽ�*<e,4���?wɽ�*<eɽ�*<eɽ�*<eɽ�*<e+�n�/�G/���?���V�mB��W�����D}���+H-KB�i𰱁�
���2Q�]�Q�Mɽ�*<eɽ�*<ex�\�uɽ�*<eɽ�*<eɽ�*<e{�<%5��*�B��;�d �����Җ LF�zN�����{�<%5� XdJA����Dtt�ɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�]Ӟve�`䷟����{v���)`���#�-KB�i𰿘P�6;7}o:����v�ɽ�*<eɽ�*<ex�\�uɽ�*<eɽ�*<eɽ�*<eɽ�*<e!�T9�u�P�+H�"�o�6�ꪕ�j7�po�W|9��\ʶ���1�%�^|��]`�Q�]�Q�Mɽ�*<eɽ�*<eNM{9q��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��r���
�JP$����Җ LF�zN�����{�<%5��g� ���Mh�]=Q�]�Q�Mɽ�*<eɽ�*<eҝ[��R�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�e��\ȟ)�;C�Q���Җ LF,ҌyX�� �ה���T�����)y���:��`ɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<eɽ�*<e�W7P�%����o=jG�7�7�Uz� �[��I�D�J�;�e(<�KB��7�1���w$o����� Fx�ɽ�*<eɽ�*<e,4���?wɽ�*<eɽ�*<eɽ�*<eɽ�*<e+�n�/�G/���?���V�mB��W�����D}���+H
j�����@��M��^��l�ɽ�*<eɽ�*<ex�\�uɽ�*<eɽ�*<eɽ�*<e��D�M��~:��#��;�d �� �ϵ%[��6ҷ�׸�م|���A6��l��1�k�ɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����^��mߠ�]�:.H.�4��vA�my�+T��u0�/���>;�# m	�ɽ�*<eɽ�*<e�VJUT���?�(<��ɽ�*<eɽ�*<e�W7P�%T��82�9��%�>v;��V�mB���x��{Ж��ٿEE)�dC��)�Ζ�ۺɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<eɽ�*<eɽ�*<eɽ�*<eșQ�z�~�AA��A�Y�sʶ��6LTy_2~��	�+T��u0���8���8��8ɽ�*<eɽ�*<e�VJUT���?�(<��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eD���p �W(�$ɯ*���S���)��Y7W��*�T��82�9!&���S+zW-;�+j8ɽ�*<eɽ�*<e����n��rɽ�*<eɽ�*<eɽ�*<eɽ�*<e��vVK�`^|��]`��V�mB���x��{Ж��ٿEE)�dC���_�av"	;��%���ɽ�*<eɽ�*<ex�\�uɽ�*<eɽ�*<eɽ�*<eɽ�*<e�2R&�N5ݐ�Mh�]=BQ��F�-�zN�������N&d�U��j��Eh����
lD��#��u��^1�������~���=���K��rq��& *R�yp��M�{�Z����q|���N\ZAܸ���R���7dj�7Y�I\���ֻ'r�f�'��Sb�&9�ΘQ�z�N̨ <�t-*�m`�| �;�e(<�KB\���ֻ'r�f�'��Sb�&9�����ڎXJ��&�+{����W&[�6���d�����8�:���2�i;�j��Eh_����nc���a5��O)ɠo>f\���ֻ'r�f�'��Sb�&9�Ο�Q5��;�D�Lw��=�zN�������N&d�U��j��Eh����
lD��#��u��^1�������~���=���Kɕ?kV7�2x!W`�lM�{�Z����q|���mVW��c�=�ﭞf��Q�Lj}���J�<A�]8��F�t�e�&�W�Lƍi�&���㗟��<�Em`�| �;�e(<�KB\���ֻ'r�f�'��Sb�&9�����ڎXJ��&�+{����W&[��E��O�-����7H���2�i;�j��Eh����
l�p������HN�E�����#4�j��Eh_����nc��E��whFo+�SZu&ꬶ�R�E�HP8jΗCf�|�D��}L�7���&S�> �1J�`���'t,�|�h�qBK�,����������n��r\���ֻ'r�f�'��Sb�&9�Ο�Q5��;B��焷sm�j��Eh_����nc���a5��m`�| �� ����o\���ֻ'r�f�'��Sb�&9�����ڎXJ��&�+{����W&[�a� ��^*��;LA��2�i;�j��Eh����
l�p����������J��%O�w`�!\���ֻ'��\yJ�	^^D�g�$�W��#T���>�K�Rɽ�*<e���J��Br(�&G!1���s�D�<@m̞���&m(��ϑi���8xH��N�ƣ��T�O�]t��j���F�t�e�&�W�Lƍ���b��{��%e�܉������F�t�e�Q��8��y	�[�xGY;�=��O��b2�M/��Jm`�| �ɽ�*<e\���ֻ'r�f�'��Sb�&9�����ڎXJ��&�+{����W&[��c�p�@L�ɽ�*<e��2�i;�j��Eh����
l�p������W�*��|��z8�2���q|���N\ZAܸ�ˀ����lv�zN�������N&d�U��j��Eh����
lD��#��u��^1�������~���=���K�[m3Eo��VJUT���M�{�Z����q|���mVW��c�=j0 �M�hh�J�.�~\���ֻ'��\yJ�	��{���b*�Nf�TJ1r���� hy������~�G:fGv���&�;���*������
nP
,����c��c�~Vp�^|��]`�չ������J��Br(�&G!1���s�D�|�u�$2�B�$D����pQcΗCf�|���G8�V���l�06��1	��S��`���%�;�+�3�q�w��ΗCf�|�D��}L�7���&S�> �1J�`���'t,�|�J���8�p��˾�[(���d֨\���ֻ'r�f�'��Sb�&9�� kdt]��8w_�}�X"n����pQcΗCf�|���G8�V�����,(Q'�!Y������� hyW|9��\�2���K,v����W���P�6;7}x`һaB�ɽ�*<eɽ�*<eɽ�*<e,4���?wdFK��/��J��oj��˩$fMT�Ҁ��O)ɠo>f��7�1��kC����k�)�Z�D�Lw��=�zN�����1稆���%A�O�����`�f ��{I����!�O1�p<�gɽ�*<eɽ�*<eɽ�*<e�VJUT���`Zʤ|�ev��</�Sb�&9�ΘQ�z�N̨ <�t-*�5��)ϋ�2���K,Ah�@�;�o��R���7<���^Z�����Ť2��9�|2���K,v����W�������h����&��ɽ�*<eɽ�*<eɽ�*<e,4���?wdFK����f0%ڡU���)ݝk,�IM�+�I����p�A�O�����D��}L�8��݌��?ɕ?kV7�hFo+�SZu�L�@�~�>�م|���T�����)�堒�c���
��R'ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r��7�1��kC����=gx�s8�8<������7�1�;��`�:މ[�xGY;����8��,*�0�ia�Y�"WoQ��;ys2Ad ݰm�H ��E��6��W��#T�m�2��&�ɽ�*<eɽ�*<eɽ�*<e[���g�Q����o=$W.����| gl�n�!�/��vJ�k�%:��</�Sb�&9��jVYFM�����>W�_��y�ճ���W7P�%����o=$W.����|�z ��>ԴW�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M,J����2���K,Ah�@�;�o�z �wB�dFK��/��J��oj��˩$fMT�Ҁ��m`�| �ɽ�*<e��7�1��kC����J��!㣝˻�%e�܉�z�iU�}ɽ�*<eɽ�*<eɽ�*<e|�'B���A�O�����D��}L�8��݌��?/���?��0�ۧ��5�dFK����f0%ڡ,��j��z�IYLy�͵�R}�&ꬶ�RQ�1	�|T�����)�堒�c�3�R�3�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r��7�1��kC�������f�άe[;Zl�fA�O�����D��}L�8��݌��?;L�?�j7ߔ��� hyW|9��\�2���K,v����W�!&���S+۳�EwW�ɽ�*<eɽ�*<eɽ�*<e,4���?wdFK����f0%ڡQ�Y�<B�$D�#�6KF5���h�!1���s�D�|�u�$2���;=6
��y�ճ���W7P�%����o=$W.����|̃��h�&,m�2��&�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M,J����2���K,Ah�@�;�o�m�[��k�%:��</�Sb�&9��f���ڳ�x�G#�S�t	�g!���Q��;ys2Ad ݰm�H ��E��6�J�EL�cm��h�n�gɽ�*<eɽ�*<eɽ�*<e[���g�Q����o=$W.����|��`��)�:/6�W��k�%:��</�Sb�&9�� kdt]��8���T�JX[��y�ճ���W7P�%����o=$W.����|�TErǃ++��c��W�����ɽ�*<eɽ�*<eɽ�*<e�M,J����2���K,6r�?x��}x���Q�0�ۧ��5�dFK����f0%ڡZm��B�R&�[��%q�5�쒈��eҥŖqW|9��\�2���K,ݥ D���z}x���Q���6�Geɽ�*<eɽ�*<eɽ�*<e,4���?wdFK����f0%ڡ)��m�SD+�?M�2D�5�O�A�O�����Sd�~�fTP�d����8�ꜟ�A��y�ճ���W7P�%����o=$W.����|�TErǃ+�\�r+�=��W�����ɽ�*<eɽ�*<eɽ�*<e�M,J����2���K,`E���փ<x@y�07Qd!p*�~��#�6KF5T�����)��� @_u}ÙEǛ'�ۄ��\��tZ�����Ť2��9�|2���K,ݥ D���z}x���Q������d<�8��ЎK�ɽ�*<eɽ�*<e,4���?wdFK����f0%ڡ)��m��R�a�G��̸B������;���}��N?�{�/z���"o��D(��Gt�em�B���&��r>�ɽ�*<edFK����f0%ڡШ6�E���f�M�
V8��+ Z�W�����ɽ�*<eɽ�*<e�:��MC�ِ�}��N�M
��iͮ���P�V?8����		%Ju9���dFK����f0%ڡZm��B�W$�.:�����<���^Q�D@�ɽ�*<e��D�MAd ݰm�Haa24�2G7���7R��ɽ�*<eɽ�*<eɽ�*<e[���g�Q����o=$W.����|�o�K��o�/�����E�����G8����o=$W.����|_�_�>_PK�`v�ZP��3_y�|�Mn�_LHwې�}��N?�{�/z���"o��D�2nq�Ř�x`һaB�ɽ�*<eɽ�*<eɽ�*<e��@�7�*T�����)�8���繬d��d��t�T�,G�k�%:Ad ݰm�H$���W 5��;�Y��##m`�| �ɽ�*<e��7�1��kC����m�@�-�F��9�:~����7X��q�ɽ�*<eɽ�*<eɽ�*<e|�'B���A�O������ʾ��
���B�F�+ ����7�1��kC����m�@�-�F�K�@V�sۄ��\��tZ�����Ť2��9�|2���K,`E���փ<�~v3�����'����V8��+ Z�W�����ɽ�*<e,4���?wdFK����f0%ڡZm��B��x��kNL������d<�Ju9���dFK����f0%ڡ� ��`Rzǅ؊��SV8��+ Zm`�| �ɽ�*<e��7�1��kC����m�@�-�F��I�|�ЮH���<���^�� �R��;ɽ�*<eɽ�*<e|�'B���A�O�����Sd�~�fTP�d����tseQ,�ٰ���˫�#�6KF5T�����)��� @_u}�r�=_V8��+ Zm`�| �ɽ�*<e�H'b6]��X�Y6����F��X
ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��~sj@�.�k�:1[��Ur�JF�k�%:Ad ݰm�H�����1�v�5�쒈�R���%�^����<�e�/����ȁă�6�Geɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w�Q�'Ws�t���>*�2D�5�O�A�O�����-�{�0Bh�{"���S����Z �jv�5�=Ď����f��6a�s��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��@�7�*T�����)C<ɓ�|*XS5�8x�XY�Q�'Ws�t:��ʵ�~e�Ʒ2�v�!w���y��h}���.�����UF:��Ҟ�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����">��f��#�C���g�@P����H�����}��N�M
��iͮ�hc�V�*��Pfɽ�*<e�i�o���tj me�S�!�(I켚<dz�Uiɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����">��f��#�C�L�PlC�V8��+ Z5��)ϋ�2���K,�"��Ѕ"�#F��8S�B���@%����Z �jv�5�=Ď����f����v��{8��ЎK�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�1��~!���T�ө���<���^���;���}��N�M
��iͮO0�-x$�nS�B���@%�܃$���)`���#�-KB�i�`�f ��{�f>;�݃۳�EwW�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ص�Y�~�R#��Sb�&9�Ο�Q5��;���-5�M|�	R��-L�kC����k�)�Z�D�Lw��=�zN�����1稆���%ҫ�0�7�v����W���R���7m��{�2�ɽ�*<eɽ�*<eɽ�*<e�VJUT���e��qb��b>�%��D2j��˩$\��М}��(H��u�6�������jU�.&��MS?�)M�L>�;>c���8�ɽ�*<e���'fLSx=��/�ч�t}�,�IM�+�In�C���2ɽ�*<eɽ�*<eɽ�*<e[���g�Q�F{N.J�M
��iͮE�����ӫo����������>�%��D2j��˩$��}��OI�BDw��?p��y�ճ���Y7W��*��F{N.J?�{�/z��s��Ɩ���7H�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M,J����!��QE�������Cw��\��������Y�~�R#��Sb�&9�ΰ��w�]�\\�����v2_�wW|9��\�!��QE���堒�c����g�#w#�o�Oɽ�*<eɽ�*<eɽ�*<e,4���?w|�	R��-L�kC����pr�΅�0ǵ�bhF_������Y�~�R#��Sb�&9��jVYFM�����>W�_��y�ճ���W7P�%�F{N.J?�{�/z�q�o�y�#ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M,J����!��QE�������C��SA>�1����{�}f�����.���p����o��@(}����ZЖ��ٿE-KB�i�`�f ��{�f>;�݃�R	V��v�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ص�Y�~�R#��Sb�&9�Ο�Q5��;��%e�܉8�̣*���-KB�i���/�T�f>;�݃f�Ӗ�F>��y�ճ���W7P�%�F{N.J?�{�/z��ȵ��,ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M,J����!��QE�������C�s�Z���ܷ��{�}f�����.���p�������/�W�܃$���)`���#�-KB�i�`�f ��{Ȯ�^q.J1����8�:�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ص�jU�.&��MS?�)^|��]`�5��)ϋ�SS���u�!1���s�D�|�u�$2���;=6
��y�ճ���W7P�%�F{N.J?�{�/z�k���CдW�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M,J����!��QE�������C��ye�|�	R��-L;��`�:މ[�xGY;�q����d�m`�| ����&�<���{�}f$W.����|Y�<d�2!#��&��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e|�'B���ҫ�0�7�Ah�@�;�o��D�\å��Bi��t�F{N.JIK�vv��8k�>�x��D�\åǓ�Lb�&ꬶ�R{�<%5��jU�.Z�?�v&i5�m�3'k:�5��;#tMɽ�*<eɽ�*<eɽ�*<e����n��r���{�}f$W.����|ar�A�D��+��c�5��)ϋ�!��QE���8����竁�F�k	�`v�ZP��3_y�|�Mn�_LHw�-KB�i�Sd�~�fT ��w����S�P'qɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ص�jU�.$���W 5�%�u�){K=�n\��{J-KB�i�Sd�~�fTP�d����8�ꜟ�A��y�ճ���W7P�%�F{N.J?�{�/z����P�V?f�,1+��+ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M,J����!��QE���8����竁�F�k	�.���Ȁ�������Sx=��/)��m�.8��l�Ʒ2�v�ɽ�*<e���'fLSx=��/Ш6�E��R�a�G��̸B��ຐ �R��;ɽ�*<eɽ�*<e[���g�Q�F{N.J�M
��iͮ���P�V?� �^J��ٰ���˫�������jU�.aa24얭�@�W������d<�xg��r��*�zN�����1稆���%ҫ�0�7�ݥ D���z}x���Q�˃�6��Rb�<dz�Uiɽ�*<eɽ�*<e�VJUT���e��qb��bSx=��/)��m���f�M�
V8��+ Z5��)ϋ�!��QE���8����竁�F�k	�"vЅ\�p;kwֹZ�����Ť2��9�|!��QE���8�����w�=*~���|��.ɽ�*<eɽ�*<eɽ�*<e,4���?w|�	R��-L�kC����m�@�-�F���{��cZy�ʏY�u�����{�}f$W.����|_�_�>_PK�`v�ZP��3_y�|�Mn�_LHw�-KB�i�Sd�~�fT^�0��ş��l�G�䗴W�����ɽ�*<eɽ�*<eɽ�*<e�����ص�jU�.aa24�ףr<$�.K-��}%��|�	R��-L�kC����pyM��]�|͈��T�<����ZЖ��ٿE-KB�i�Sd�~�fT^�0��şAwo��o�Aв�2Gɽ�*<eɽ�*<eɽ�*<e�����ص�jU�.$���W 5��I>/�4	�!�L?7Ƌҫ�0�7�`E���փ<�v�F�
o��U�����m`�| �ɽ�*<e���{�}f$W.����|�o�K��o��������!�(I켚<dz�Uiɽ�*<eɽ�*<e|�'B���ҫ�0�7�`E���փ<�v�F�
o���'����V8��+ Z5��)ϋ�!��QE����� @_u}c�XO�_ag�̸B���Q�D@�ɽ�*<e���'fLSx=��/Zm��B��H�@�p1˃�6��Rb�<dz�Uiɽ�*<eɽ�*<e[���g�Q�F{N.J?�{�/z���"o��DI>5}�%@lV8��+ Z5��)ϋ�!��QE����� @_u}�r�=_V8��+ Zm`�| �ɽ�*<e�H'b6]�i��m�O�!f�� �fɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��~sj@	c�W.�ҽl��P�ti+8�̣*���-KB�i�-�{�0B'��U0D9h��b���c��Gj�B��{���	��8��㵒���8�:�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e!��$и3��/�Ѭ�}��&�rS5��)ϋ�!��QE��C<ɓ�|*X�i��g��Z�������0{�I�/�ʸ�}4Wj̼��Aв�2Gɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w|�	R��-L�kC����d5K�;���2y�H�1�ϱ���V#�E:~�9�[�P9��7�r��s�ݚ}� .=2�����g�@P�M�tb�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�H'b6]R�U�(�N,�o��v������jU�..���~�$�6��V^�����Z �jv�5�=�1�ϱ�d� �c�#�!�(I켚<dz�Uiɽ�*<eɽ�*<eɽ�*<eɽ�*<e�1��~!ځ�Ex���L�PlC�V8��+ Z5��)ϋ�!��QE��C<ɓ�|*X�����d<�xg��r��*�zN������%,!u�r�	c�W.�ҽ��*�jCe�V8��+ Z�W�����ɽ�*<eɽ�*<eɽ�*<e�VJUT���Օ�^�e�{��������v��{Ju9���|�	R��-L�kC����}PYg��?V8��+ Zm`�| �;�e(<�KBIή�%`��kC����J��!㣝˰T�+Tnɽ�*<eɽ�*<eɽ�*<eɽ�*<e|�'B���)�ߙmit�D��}L�8��݌��?/���?��5��)ϋ�}%^Y[�\VAh�@�;�o��P�6;7}z�s]eNN`ɽ�*<edFK��Z
�i(�?;~�)�D?R��9����h�n�gɽ�*<eɽ�*<eɽ�*<e�:��MC��
j���IK�vv��8k�>�x��R���7dj�7Y�IIή�%`��kC�������K�@w� <�t-*�m`�| �ɽ�*<eIή�%`��kC�����Έx�3�㗟��<�E�W�����ɽ�*<eɽ�*<eɽ�*<e|�'B���)�ߙmit����/�T�>��܎�^�7a0b�dFK���e�: z�[j��˩$��}��OI�BDw��?p��y�ճ���Y7W��*������x�$W.����|txG�z��h�CÁ�� ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M,J����}%^Y[�\VAh�@�;�o���
���25��)ϋ�}%^Y[�\VmVW��c�=3��,�����] �, ����Z~�0�V�a
j���?�{�/z�wM�.����*��;LAɽ�*<eɽ�*<eɽ�*<eɽ�*<e��@�7�*�-H嵰. �����C���g�#wf��h�\
j���IK�vv��8k�>�x�Д�٪,�j�M��gt&ꬶ�RQ�1	�|�-H嵰. �堒�c�}�/͓ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rIή�%`��kC����k�)�Z!�"
��u)�ߙmit�D��}L�8��݌��?°�:_��Z�����Ť2��9�|}%^Y[�\Vv����W���P�6;7}��H�8�ɽ�*<eɽ�*<eɽ�*<e,4���?wdFK���e�: z�[j��˩$fMT�Ҁ����T�O�!�"
��u)�ߙmit����/�T�f>;�݃f�Ӗ�F>��y�ճ���W7P�%�����x�$W.����|���p�w��W�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M,J����}%^Y[�\VAh�@�;�o�a7���\dFK���e�: z�[j��˩$&6��u48m`�| �;�e(<�KBIή�%`��kC�����z��=��3��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e|�'B���)�ߙmit����/�TȮ�^q.J1Ը�x-L
������x������.���p�����l�06��1	��S��`&ꬶ�RQ�1	�|�-H嵰. �堒�c��[m3Eo�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rIή�%`��kC����(� ��ڷ4-V�]�+ٯ
j���IK�vv��8k�>�x�}IU��	����Zq1Q�e
j���?�{�/z��QT�G$aW��)f�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��@�7�*�-H嵰. �����C�[�eonD�Ƣ2�S�
j���IK�vv��8k�>�x��D�\åǓ�Lb�&ꬶ�RQ�1	�|�-H嵰. yyֶ�T@�����n����z#U�9�ɽ�*<eɽ�*<eɽ�*<e����n��rIή�%`��kC�����V�j�Mc(J ��!�"
��u)�ߙmit��Sd�~�fTP�d�����M`.�m`�| ���{c^��Iή�%`��kC����K��H7E������W�����ɽ�*<eɽ�*<eɽ�*<e|�'B���)�ߙmit���ʾ�� ��w���-��}%��dFK��Z
�i(�?Zm��B�'y!~ޓ�m1	��S��`&ꬶ�RQ�1	�|�-H嵰. yyֶ�T@ÙEǛ'��7X��q�ɽ�*<eɽ�*<eɽ�*<e����n��rIή�%`��kC����m�@�-�F��qA�KJ���
�,��,�����x�$W.����|ar�A�D���\�r+�=�m`�| �ɽ�*<eIή�%`��kC����K��H7Z�j"�nm�B����h�n�gɽ�*<eɽ�*<e|�'B���)�ߙmit���ʾ�� ��w���"�#F��8k�kN�$߈k�%:A�^_p�xaa24얭�@�W������d<�xg��r��*�zN�����1稆���%)�ߙmit��Sd�~�fT ��w����"vЅ\�����}g�ɽ�*<eɽ�*<e�VJUT���`Zʤ|�evA�^_p�x$���W 5�~��/��K�am@���H�(�)�ߙmit��Sd�~�fTP�d�������q�ޤS�B���@%����ZЖ��ٿE
j���?�{�/z���"o��D�$@�՛��z�iU�}ɽ�*<eɽ�*<eɽ�*<e��@�7�*�-H嵰. �8���繬d��d�2���m�#�6KF5�-H嵰. ��� @_u}}!�Lڜ<��q��M�"���tI�tQ��;ys2A�^_p�xaa24�2G7����S�P'qɽ�*<eɽ�*<eɽ�*<e[���g�Q�����x�$W.����|�o�K��o�����ﴖ=�n\��{J
j����M
��iͮ�5�MP���i��g��Z�����Ť2��9�|}%^Y[�\V`E���փ<�~v3����U������W�����ɽ�*<eɽ�*<e,4���?wdFK��Z
�i(�?� ��`RzǍ�����5��)ϋ�}%^Y[�\V`E���փ<�v�F�
o��U�����m`�| �ɽ�*<eIή�%`��kC����m�@�-�F�4�)�*�z�G5�td'����}g�ɽ�*<eɽ�*<e|�'B���)�ߙmit��Sd�~�fTP�d����{M�y0��bm�B�����H�(�)�ߙmit���ʾ�֓��P2��G5�td'p;kwֹZ�����Ť2��9�|}%^Y[�\V`E���փ<�~v3��G������r��5p���ɽ�*<eɽ�*<e,4���?wdFK��Z
�i(�?Zm��B��x��kNL�˃�6��Rb8�>��z������x�$W.����|_�_�>_PK�"vЅ\�p;kwֹZ�������0{�I�S�B���k��X�Y6����F��X
ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w�Q�'Ws�t�0�]`~WF[��Ur�JF�k�%:A�^_p�x�����1�v�5�쒈�R���%�^����<�e�/�S�B���k}��&�rS�W�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w�Q�'Ws�t�0�]`~WF-��}%��dFK��Z
�i(�?�l8�Բ��� �ɽ�*<e�i�o��� PزK`Q�6a�s��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e[���g�Q�����x�$W.����|+�<b�g�fq�ٓ @ӱ��n�:��ʵ�~e�Ʒ2�v�!w���y��h}��� PزK`Q[���MĞ�>υU�%ߏɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����">�{���	��=���n���jX.�k�%:A�^_p�x.���~�$�6��V^�����Z �jv�5�=�1�ϱ�a�9�5���!�(I켚<dz�Uiɽ�*<eɽ�*<eɽ�*<eɽ�*<e�1��~!���MY���L�PlC�V8��+ Z5��)ϋ�}%^Y[�\V�"��Ѕ"�#F��8S�B���@%����Z �jv�5�=�1�ϱ�-ڲ�TrM��K�am@���h�n�gɽ�*<eɽ�*<eɽ�*<eɽ�*<e�1��~!���MY�ޡ�W���k�kN�$߈k�%:A�^_p�xT����=����<���^Q�D@��g����j�1���,S��c�P2� ����N�`?=ɽ�*<eɽ�*<eɽ�*<eɽ�*<e[���g�Q7��ɇ�F������.���p����y�P����g=�n\��{J8�|q{+��M
��iͮeg�/�1	��S��`&ꬶ�RxP�Z�W揉ry�k��堒�c���rq��&�:8[�d�-ɽ�*<eɽ�*<eɽ�*<e����n��rn�>�B";��`�:މ[�xGY;�ZQ�R�"=����+�GB��,d�?��S��c�P&��MS?�)M�L>�;>c���8�ɽ�*<e�@����S��c�P94���i�Lj}�����7H�ɽ�*<eɽ�*<eɽ�*<e[���g�Q7��ɇ�F�$W.����|�rR��`~�:���y��VX�
�j�3�)򢦃�v!1���s�DC��ŀ�~,�IM�+�I�$�l� ��2]|B�~W��Z0B��)�xoĪ���D�	�Ӯ#�3"�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�:��MC��8�|q{+��M
��iͮ�s��ƖO�bJŤ<�8�|q{+�IK�vv��8k�>�x���
���2m`�| �� ����on�>�B"�kC�����ݮ5q.u�[0��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e|�'B������H��6���/�T`xr�a�%O�w`�!n�>�B";��`�:މ[�xGY;�V�3yn�3����m�c�zN�����1稆���%���H��6`�f ��{�Hb�0"	ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT������9f?S��c�PD!�yk��	vO���S7��ɇ�F������.���p����o��@(}����ZЖ��ٿE8�|q{+�?�{�/z�eg�/�b2�M/��J�W�����ɽ�*<eɽ�*<eɽ�*<e�iƅ��)򢦃�v!1���s�D�׸ǭ��?��z�IYLy����G87��ɇ�F�$W.����|Tu������T�O���ʶ��^�ɽ�*<e��Z0B��)�xoĪ��8�z4�����iuɽ�*<eɽ�*<eɽ�*<eɽ�*<e�:��MC��8�|q{+��M
��iͮ6s��}�X�
�j�3�)򢦃�v!1���s�D<��M�D����V��g����j�1���,S��c�PL����^|��]`�W�����ɽ�*<eɽ�*<eɽ�*<e[���g�Q7��ɇ�F�$W.����|�E��Cӽ��}Mxw��Z0B������3�j��˩$�ܚ����t)��`�zN�����1稆���%���H��6`�f ��{o�Wq�AGɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT������9f?S��c�P&��MS?�)hh�J�.�~n�>�B";��`�:މ[�xGY;�q����d�m`�| ����&�<n�>�B"�kC�����o�2��vc �?Y*ɽ�*<eɽ�*<eɽ�*<eɽ�*<e|�'B������H��6���/�T�A�c���렗k"f+n�>�B";��`�:މ[�xGY;���e�8��������d�zN�����1稆���%���H��6�Sd�~�fT ��w���7R��ɽ�*<eɽ�*<eɽ�*<e�VJUT������9f?S��c�P$���W 5�m�3'k:�����G87��ɇ�F�$W.����|�o�K��o��rK-�'��<��q��M�"���tI�tj�1���,S��c�PZ�?�v&i5%�u�){K۳�EwW�ɽ�*<eɽ�*<eɽ�*<e[���g�Q7��ɇ�F�$W.����|ar�A�D��^ţ�U�X�
�j�3�ry�k��8����竁�F�k	�{d��T��zN�����1稆���%���H��6�Sd�~�fT ��w���b:n\��ɽ�*<eɽ�*<eɽ�*<e�VJUT������9f?S��c�Paa24얭�@�W�S5�8x�XY��Z0B��)�xoĪ)��m�.8��l�Ʒ2�v�ɽ�*<e�@����S��c�PZ�?�v&i5Pn���&���!�(I켚<dz�Uiɽ�*<eɽ�*<e[���g�Q7��ɇ�F�$W.����|ar�A�D��3��|��V8��+ Z5��)ϋ��z��X3�`E���փ<x@y�07Q���:��e
���4�Qp?��y�ճ���W7P�%7��ɇ�F�$W.����|�TErǃ+����%֎�5p���ɽ�*<eɽ�*<eɽ�*<e�M,J���܇z��X3�6r�?x��}x���Q�˃�6��Rb8�>��z�7��ɇ�F�$W.����|�o�K��o�E���@��V8��+ Zm`�| �ɽ�*<en�>�B"�kC����m�@�-�F�]��?�`C���z#U�9�ɽ�*<eɽ�*<eɽ�*<e|�'B������H��6�Sd�~�fTP�d����91��?��!�"
��u���H��6��ʾ��B`�M�5�쒈��eҥŖqW|9��\ʇz��X3�`E���փ<�~v3��`@T�;�/ɽ�*<eɽ�*<eɽ�*<e,4���?w��Z0B��)�xoĪZm��B��x��kNL�O)ɠo>fn�>�B"�kC����pyM��]�|͈��T�<����ZЖ��ٿE8�|q{+�?�{�/z���"o��D��Q(�>·�ۃRIɽ�*<eɽ�*<eɽ�*<e�iƅ��ry�k���� @_u}�z�`u�t�,��/8�|q{+�?�{�/z���"o��D/��	���Ʒ2�v�ɽ�*<e�@����S��c�Paa24�2G7���"�#F��8��5p���ɽ�*<eɽ�*<e[���g�Q7��ɇ�F�$W.����|�o�K��o�<�3�N��!�(I�8�>��z�7��ɇ�F�$W.����|_�_�>_PK"�#F��8S�B���@%����ZЖ��ٿE8�|q{+�?�{�/z���"o��D�Z�9�V8��+ Z�W�����ɽ�*<eɽ�*<e�iƅ��ry�k��8���繬d��d��V��P ��Ju9�����Z0B��)�xoĪ� ��`Rz�6vZ�%�MS�B���@%����Z �jv�5�=�1�ϱ��9j�`�<R5��;#tMɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�1��~!hsrTq�m��~-y75��)ϋ��z��X3��"��Ѕ�`v�ZP��3_y�|��K[+��1�ϱ�1m e�۳�EwW�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�1��~!hsrTq�m�����7X�
�j�3�ry�k�C<ɓ�|*X�i��g��Z�������0{�I����d�J4Wj̼��Aв�2Gɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��Z0B��)�xoĪ��eo6����ɒ(�{���	����	Y�[�ۄ��\��t\���OxO���<�e�/����d�J2�����j�m���[̹ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w�Q�'Ws�t'�'�N��q��K�`5��)ϋ��z��X3��"��Ѕ��K�`m`�| �ɽ�*<e�H'b6]~s>B`LjP�����d<�8��ЎK�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��~sj@�c��y�-��Mbg(�!�̸B������;��8�|q{+��M
��iͮf��}J!W-V8��+ Zm`�| �ɽ�*<e�H'b6]~s>B`LjP˃�6��Rb�<dz�Uiɽ�*<eɽ�*<eɽ�*<eɽ�*<e��~sj@�c��y�-�J\O�Z�V8��+ Z5��)ϋ��z��X3��"��Ѕ�"vЅ\�p;kwֹ���� hyW|9��\ʁ����=�v����W���P�6;7}x`һaB�ɽ�*<eɽ�*<eɽ�*<e,4���?w��Z0B��381�Mj��˩$fMT�Ҁ��O)ɠo>f|2w�e�Q��kC����k�)�Z�D�Lw��=�zN�����1稆���%�I�\�m��`�f ��{I����!�O1�p<�gɽ�*<eɽ�*<eɽ�*<e�VJUT������9f?Q90y0�ȐSb�&9�ΘQ�z�N̨ <�t-*�5��)ϋ������=�Ah�@�;�o��R���7<���^Z�����Ť2��9�|�����=�v����W�������h����&��ɽ�*<eɽ�*<eɽ�*<e,4���?w��Z0B������?U���)ݝk,�IM�+�I����p��I�\�m��D��}L�8��݌��?ɕ?kV7�hFo+�SZu�L�@�~�>aV�CF�[^��,Fwp�堒�c���
��R'ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r|2w�e�Q��kC����=gx�s8�8<����|2w�e�Q�;��`�:މ[�xGY;����8��,*�0�ia�Y�"Woj�1���,���Lt�c� ��E��6��W��#T�m�2��&�ɽ�*<eɽ�*<eɽ�*<e[���g�QRIꐦO�j$W.����| gl�n�!�/��vJ��,d�?��Q90y0�ȐSb�&9��jVYFM�����>W�_��y�ճ���W7P�%RIꐦO�j$W.����|�z ��>ԴW�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M,J���܁����=�Ah�@�;�o�z �wB���Z0B��381�Mj��˩$fMT�Ҁ��m`�| �ɽ�*<e|2w�e�Q��kC����J��!㣝˻�%e�܉�z�iU�}ɽ�*<eɽ�*<eɽ�*<e|�'B����I�\�m��D��}L�8��݌��?/���?��0�ۧ��5���Z0B������?,��j��z�IYLy�͵�R}�&ꬶ�RxP�Z�W�^��,Fwp�堒�c�3�R�3�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r|2w�e�Q��kC�������f�άe[;Zl�f�I�\�m��D��}L�8��݌��?;L�?�j7ߔ��� hyW|9��\ʁ����=�v����W�!&���S+۳�EwW�ɽ�*<eɽ�*<eɽ�*<e,4���?w��Z0B������?Q�Y�<B�$DX�
�j�39��#l��B!1���s�D�|�u�$2���;=6
��y�ճ���W7P�%RIꐦO�j$W.����|̃��h�&,m�2��&�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M,J���܁����=�Ah�@�;�o�m�[���,d�?��Q90y0�ȐSb�&9��f���ڳ�x�G#�S�t	�g!���j�1���,���Lt�c� ��E��6�J�EL�cm��h�n�gɽ�*<eɽ�*<eɽ�*<e[���g�QRIꐦO�j$W.����|��`��)�:/6�W���,d�?��Q90y0�ȐSb�&9�� kdt]��8���T�JX[��y�ճ���W7P�%RIꐦO�j$W.����|�TErǃ++��c��W�����ɽ�*<eɽ�*<eɽ�*<e�M,J���܁����=�6r�?x��}x���Q�0�ۧ��5���Z0B������?Zm��B�R&�[��%q�5�쒈��eҥŖqW|9��\ʁ����=�ݥ D���z}x���Q���6�Geɽ�*<eɽ�*<eɽ�*<e,4���?w��Z0B������?)��m�SD+�?M�2D�5�O��I�\�m�ʹSd�~�fTP�d����8�ꜟ�A��y�ճ���W7P�%RIꐦO�j$W.����|�TErǃ+�\�r+�=��W�����ɽ�*<eɽ�*<eɽ�*<e�M,J���܁����=�`E���փ<x@y�07Qd!p*�~�X�
�j�3^��,Fwp��� @_u}ÙEǛ'�ۄ��\��tZ�����Ť2��9�|�����=�ݥ D���z}x���Q������d<�8��ЎK�ɽ�*<eɽ�*<e,4���?w��Z0B������?)��m��R�a�G��̸B������;���	�d�?�{�/z���"o��D(��Gt�em�B���&��r>�ɽ�*<e��Z0B������?Ш6�E���f�M�
V8��+ Z�W�����ɽ�*<eɽ�*<e�:��MC�ِ�	�d��M
��iͮ���P�V?8����		%Ju9�����Z0B������?Zm��B�W$�.:�����<���^Q�D@�ɽ�*<e�@�������Lt�c�aa24�2G7���7R��ɽ�*<eɽ�*<eɽ�*<e[���g�QRIꐦO�j$W.����|�o�K��o�/�����E�����G8RIꐦO�j$W.����|_�_�>_PK�`v�ZP��3_y�|�Mn�_LHwې�	�d�?�{�/z���"o��D�2nq�Ř�x`һaB�ɽ�*<eɽ�*<eɽ�*<e�iƅ�^��,Fwp�8���繬d��d��t�T�,G��,d�?����Lt�c�$���W 5��;�Y��##m`�| �ɽ�*<e|2w�e�Q��kC����m�@�-�F��9�:~����7X��q�ɽ�*<eɽ�*<eɽ�*<e|�'B����I�\�m�ʽ�ʾ��
���B�F�+ ��|2w�e�Q��kC����m�@�-�F�K�@V�sۄ��\��tZ�����Ť2��9�|�����=�`E���փ<�~v3�����'����V8��+ Z�W�����ɽ�*<e,4���?w��Z0B������?Zm��B��x��kNL������d<�Ju9�����Z0B������?� ��`Rzǅ؊��SV8��+ Zm`�| �ɽ�*<e|2w�e�Q��kC����m�@�-�F��I�|�ЮH���<���^�� �R��;ɽ�*<eɽ�*<e|�'B����I�\�m�ʹSd�~�fTP�d����tseQ,�ٰ���˫�X�
�j�3^��,Fwp��� @_u}�r�=_V8��+ Zm`�| �ɽ�*<e�H'b6]��CVD�!f�� �fɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��~sj@u��^��^�l��P�ti+8�̣*��ؐ�	�d��M
��iͮ9n��5�m`�| ��C4�XȓH'b6]��CVD��6�Geɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��~sj@u��^��^����>*�2D�5�O��I�\�m�ʃ-�{�0Bh�{"���S����Z �jv�5�=�1�ϱ�D�5�1T\传]�RH�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�iƅ�^��,FwpC<ɓ�|*XS5�8x�XY�Q�'Ws�t���������P�7rV�܃$����5wz��pN�1�ϱ��I<t^8Q0:��Ҟ�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�1��~!��y��;ڽ��g�@P����H�����	�d��M
��iͮ�hc�V�*��Pfɽ�*<e�i�o����utm&Yj�s|Oݽ㺢�"��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����">�{���	��c�L�ϼ^G5�td'���ֿ74�|2w�e�Q��kC������7�we*�̸B���Q�D@�ɽ�*<e�i�o����utm&Y���v��{8��ЎK�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����">�{���	���f�&��\���<���^���;���	�d��M
��iͮO0�-x$�nS�B���@%�܃$���)`���#���Jnj��?�{�/z�eg�/�����8�:�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�iƅ����v%�|!1���s�D�׸ǭ��?�a3#L����,d�?���;�TD!�yk��c�����y�ճ���W7P�%t���̌$W.����|�.k-���!!�u�"J�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M,J����ڇ��C�mVW��c�=j0 �M�M�L>�;>cnn37��m��Jnj���M
��iͮ�&�ϔ��5�B�������ZЖ��ٿE��Jnj��?�{�/z�E�����vL���5ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�iƅ�Ɖ�D��0L�����Cɕ?kV7� 3�/
B�St���̌�����.���p�������t�i���+Ȉ4�mJ�KW�B�	E�7��+ v��`�f ��{�q�
<~�n�C���2ɽ�*<eɽ�*<eɽ�*<e�VJUT������9f?��;�TBx�Ğ��ɘ�n�e�j���,d�?���`��MǐSb�&9�ΰ��w�]�\\�����v2_�wW|9��\�ڇ��C�v����W��Д�٪,�
E�iU�)ɽ�*<eɽ�*<eɽ�*<e,4���?w��Z0B��n�Rd%�I��s�$���b\	y`�5��)ϋ�ڇ��C�mVW��c�=����E��ݼW��#T���>�K�Rɽ�*<e��Z0B��n�Rd%��K��Ɛα,������ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�:��MC�ٌ�Jnj���M
��iͮ��s<%��X�
�j�3���v%�|!1���s�D�׸ǭ��?y*����iɽ�*<e�@������;�T2� ���_d�Ǹ����z#U�9�ɽ�*<eɽ�*<eɽ�*<e[���g�Qt���̌�����.���p����y�P����g����!�X�
�j�3Ɖ�D��0L�����C/���?��bb����G�zN�����1稆���%��+ v��`�f ��{�^�WvQt�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT������9f?��;�T9v5���6���k�t���̌�����.���p�������/�W�܃$���)`���#���Jnj��?�{�/z�k���CЃ�6�Geɽ�*<eɽ�*<eɽ�*<eɽ�*<e�iƅ�Ɖ�D��0L�����Ci���!�)�2D�5�O㉾+ v��D��}L�8��݌��?i���!�)�z�s]eNN`ɽ�*<e��Z0B��n�Rd%�X�(��8
c?�4c
�}�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�:��MC�ٌ�Jnj���M
��iͮk���C�5��)ϋ�ڇ��C�mVW��c�=j0 �MފNf�TJ1rz5���W|9��\�ڇ��C�v����W���D�\å@��7�6ɽ�*<eɽ�*<eɽ�*<e,4���?w��Z0B��n�Rd%�������t���˾�[(5��)ϋ�ڇ��C�mVW��c�=����E���J�EL�cm&��r>�ɽ�*<e��Z0B��n�Rd%�Ш6�E���hƁ�,�z�iU�}ɽ�*<eɽ�*<eɽ�*<e�:��MC�ٌ�Jnj���M
��iͮ���P�V?��a��{e�X�
�j�3Ɖ�D��0L�8����竁�F�k	�`v�ZP��3_y�|�Mn�_LHwی�Jnj��?�{�/z����P�V?���Jr8�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�iƅ�Ɖ�D��0L��� @_u}E%��D�&Ը�x-L
�t���̌$W.����|�o�K��o�Z�H[�MF�z�s]eNN`ɽ�*<e��Z0B��n�Rd%�Ш6�E�.8��l·�ۃRIɽ�*<eɽ�*<eɽ�*<e�:��MC�ٌ�Jnj��?�{�/z���"o��D�>��y��!�L?7Ƌ��+ v����ʾ�� ��w���P�7rV����ZЖ��ٿE��Jnj��?�{�/z����P�V?� �^J�����"��ɽ�*<eɽ�*<eɽ�*<e�iƅ�Ɖ�D��0L��� @_u}����^EG5�td'���ֿ74�;K�Raz�kC����m�@�-�F�L�v:��!�(I�o� ���&ꬶ�RxP�Z�W�Ɖ�D��0Lyyֶ�T@��PO�K����<���^�� �R��;ɽ�*<eɽ�*<e����n��r;K�Raz�kC�����V�j��B5+o=�ٰ���˫�X�
�j�3Ɖ�D��0L�8����竁�F�k	�"vЅ\�p;kwֹZ�����Ť2��9�|ڇ��C�`E���փ<�~v3��>|
ϒ��޴W�����ɽ�*<eɽ�*<e,4���?w��Z0B��n�Rd%�Zm��B��x��kNL�0�ۧ��5���Z0B��n�Rd%�� ��`Rz�� b��m`�| ���{c^��;K�Raz�kC����m�@�-�F�^�� ���8�:�ɽ�*<eɽ�*<eɽ�*<e|�'B�����+ v���Sd�~�fTP�d���ͼ�l�G��5��)ϋ�ڇ��C�6r�?x��C'�K��w���� �ɽ�*<e�@������;�Taa24�2G7���b:n\��ɽ�*<eɽ�*<eɽ�*<e[���g�Qt���̌$W.����|_�_�>_PK�.���Ȁ���,d�?���;�Taa24�ףr<$�.K�P�7rV����ZЖ��ٿE��Jnj��?�{�/z���"o��D j��c�̸B��ຐ �R��;ɽ�*<eɽ�*<e�iƅ�Ɖ�D��0L�8���繬d��d��ym��Aٰ���˫�X�
�j�3Ɖ�D��0L��� @_u}c�XO�_ag�̸B���Q�D@�ɽ�*<e�@������;�Taa24�2G7����"vЅ\�����}g�ɽ�*<eɽ�*<e[���g�Qt���̌$W.����|�o�K��o����/*� ��K�am@���H�(𥉾+ v����ʾ�֠/��Z �^���<���^Q�D@�ɽ�*<e�i�o����_��/�d�X P��>d}ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����">�{���	��Y��y�e�ʏY�u��;K�Raz�kC����]oN�	�L�<��q��M�ZGǦ��4�h}����_��/�d˕�5_m��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����">�{���	��Z���Z��Ը�x-L
�t���̌$W.����|r3s��m`�| �ɽ�*<e�H'b6]��O0�|���QFb�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e|�'B�����+ v���-�{�0B;���7d�^����on�Q:�����.�NHm`�| ���Da�rF�H'b6]��O0�|݁��!8ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��~sj@
	}�%I^�9	��͟.O@�;K�Raz�kC����5ٗάŻV��X��xB�Z�������0{�I��IÎȌ���\�m�B����h�n�gɽ�*<eɽ�*<eɽ�*<e,4���?w�Q�'Ws�t�S���y�"�#F��8k�kN�$���,d�?���;�T���I."lkG5�td'p;kwֹZ�������0{�I��IÎ�+��%ƺ��"��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w�Q�'Ws�t�S���y��"vЅ\����ֿ74�;K�Raz�kC����}PYg��?V8��+ Zm`�| �;�e(<�KB��3����kC����J��!㣝˰T�+Tnɽ�*<eɽ�*<eɽ�*<eɽ�*<e|�'B������]-��D��}L�8��݌��?/���?��5��)ϋ�������Ah�@�;�o��P�6;7}z�s]eNN`ɽ�*<e��Z0B��N'�����;~�)�D?R��9����h�n�gɽ�*<eɽ�*<eɽ�*<e�:��MC��|m9T�g�RIK�vv��8k�>�x��R���7dj�7Y�I��3����kC�������K�@w� <�t-*�m`�| �ɽ�*<e��3����kC�����Έx�3�㗟��<�E�W�����ɽ�*<eɽ�*<eɽ�*<e|�'B������]-�����/�T�>��܎�^�7a0b���Z0B��s��g���j��˩$��}��OI�BDw��?p��y�ճ���Y7W��*��ϝO�}�$W.����|txG�z��h�CÁ�� ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M,J����������Ah�@�;�o���
���25��)ϋ�������mVW��c�=3��,�����] �, ����Z~�0�V�a|m9T�g�R?�{�/z�wM�.����*��;LAɽ�*<eɽ�*<eɽ�*<eɽ�*<e�iƅ�q>��Z�.����C���g�#wf��h�\|m9T�g�RIK�vv��8k�>�x�Д�٪,�j�M��gt&ꬶ�RxP�Z�W�q>��Z�.�堒�c�}�/͓ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r��3����kC����k�)�Z!�"
��u���]-��D��}L�8��݌��?°�:_��Z�����Ť2��9�|������v����W���P�6;7}��H�8�ɽ�*<eɽ�*<eɽ�*<e,4���?w��Z0B��s��g���j��˩$fMT�Ҁ����T�O�!�"
��u���]-�����/�T�f>;�݃f�Ӗ�F>��y�ճ���W7P�%�ϝO�}�$W.����|���p�w��W�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M,J����������Ah�@�;�o�a7���\��Z0B��s��g���j��˩$&6��u48m`�| �;�e(<�KB��3����kC�����z��=��3��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e|�'B������]-�����/�TȮ�^q.J1Ը�x-L
��ϝO�}������.���p�����l�06��1	��S��`&ꬶ�RxP�Z�W�q>��Z�.�堒�c��[m3Eo�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r��3����kC����(� ��ڷ4-V�]�+ٯ|m9T�g�RIK�vv��8k�>�x�}IU��	����Zq1Q�e|m9T�g�R?�{�/z��QT�G$aW��)f�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�iƅ�q>��Z�.����C�[�eonD�Ƣ2�S�|m9T�g�RIK�vv��8k�>�x��D�\åǓ�Lb�&ꬶ�RxP�Z�W�q>��Z�.�yyֶ�T@�����n����z#U�9�ɽ�*<eɽ�*<eɽ�*<e����n��r��3����kC�����V�j�Mc(J ��!�"
��u���]-���Sd�~�fTP�d�����M`.�m`�| ���{c^�ܖ�3����kC����K��H7E������W�����ɽ�*<eɽ�*<eɽ�*<e|�'B������]-����ʾ�� ��w���-��}%����Z0B��N'�����Zm��B�'y!~ޓ�m1	��S��`&ꬶ�RxP�Z�W�q>��Z�.�yyֶ�T@ÙEǛ'��7X��q�ɽ�*<eɽ�*<eɽ�*<e����n��r��3����kC����m�@�-�F��qA�KJ���
�,��,�ϝO�}�$W.����|ar�A�D���\�r+�=�m`�| �ɽ�*<e��3����kC����K��H7Z�j"�nm�B����h�n�gɽ�*<eɽ�*<e|�'B������]-����ʾ�� ��w���"�#F��8k�kN�$���,d�?���Ժ��h�aa24얭�@�W������d<�xg��r��*�zN�����1稆���%���]-���Sd�~�fT ��w����"vЅ\�����}g�ɽ�*<eɽ�*<e�VJUT������9f?��Ժ��h�$���W 5�~��/��K�am@���H�(𥁀�]-���Sd�~�fTP�d�������q�ޤS�B���@%����ZЖ��ٿE|m9T�g�R?�{�/z���"o��D�$@�՛��z�iU�}ɽ�*<eɽ�*<eɽ�*<e�iƅ�q>��Z�.��8���繬d��d�2���mX�
�j�3q>��Z�.���� @_u}}!�Lڜ<��q��M�"���tI�tj�1���,��Ժ��h�aa24�2G7����S�P'qɽ�*<eɽ�*<eɽ�*<e[���g�Q�ϝO�}�$W.����|�o�K��o�����ﴖ=�n\��{J|m9T�g�R�M
��iͮ�5�MP���i��g��Z�����Ť2��9�|������`E���փ<�~v3����U������W�����ɽ�*<eɽ�*<e,4���?w��Z0B��N'����ՙ ��`RzǍ�����5��)ϋ�������`E���փ<�v�F�
o��U�����m`�| �ɽ�*<e��3����kC����m�@�-�F�4�)�*�z�G5�td'����}g�ɽ�*<eɽ�*<e|�'B������]-���Sd�~�fTP�d����{M�y0��bm�B�����H�(𥁀�]-����ʾ�֓��P2��G5�td'p;kwֹZ�����Ť2��9�|������`E���փ<�~v3��G������r��5p���ɽ�*<eɽ�*<e,4���?w��Z0B��N'�����Zm��B��x��kNL�˃�6��Rb8�>��z��ϝO�}�$W.����|_�_�>_PK�"vЅ\�p;kwֹZ�������0{�Io,�)Nk���X�Y6����F��X
ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w�Q�'Ws�tC�ypVq�[��Ur�JF��,d�?���Ժ��h������1�v�5�쒈�R���%�^����<�e�/o,�)Nk�}��&�rS�W�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w�Q�'Ws�tC�ypVq�-��}%����Z0B��N'������l8�Բ��� �ɽ�*<e�i�o���lC�z�q��6a�s��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e[���g�Q�ϝO�}�$W.����|+�<b�g�fq�ٓ @�z��d��Q:��ʵ�~e�Ʒ2�v�!w���y��h}���lC�z�q�[���MĞ�>υU�%ߏɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����">�{���	���$I�-AO���jX.��,d�?���Ժ��h�.���~�$�6��V^�����Z �jv�5�=�1�ϱ�������F�!�(I켚<dz�Uiɽ�*<eɽ�*<eɽ�*<eɽ�*<e�1��~!��I;P��E�L�PlC�V8��+ Z5��)ϋ��������"��Ѕ"�#F��8S�B���@%����Z �jv�5�=�1�ϱ�ȂQ�m�K�am@���h�n�gɽ�*<eɽ�*<eɽ�*<eɽ�*<e�1��~!��I;P��E��W���k�kN�$���,d�?���Ժ��h�T����=����<���^Q�D@��g����j�1���,d������2� ����N�`?=ɽ�*<eɽ�*<eɽ�*<eɽ�*<e[���g�Q(�2Y�ǫ�����.���p����y�P����g=�n\��{J;i���`C>�M
��iͮeg�/�1	��S��`&ꬶ�RxP�Z�W揗���N�B�堒�c���rq��&�:8[�d�-ɽ�*<eɽ�*<eɽ�*<e����n��r��f�|L;��`�:މ[�xGY;�ZQ�R�"=����+�GB��,d�?��d������&��MS?�)M�L>�;>c���8�ɽ�*<e�@����d������94���i�Lj}�����7H�ɽ�*<eɽ�*<eɽ�*<e[���g�Q(�2Y�ǫ$W.����|�rR��`~�:���y��VX�
�j�3��9O�d�!1���s�DC��ŀ�~,�IM�+�I�$�l� ��2]|B�~W��Z0B�񇍞S,��m���D�	�Ӯ#�3"�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�:��MC��;i���`C>�M
��iͮ�s��ƖO�bJŤ<�;i���`C>IK�vv��8k�>�x���
���2m`�| �� ����o��f�|L�kC�����ݮ5q.u�[0��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e|�'B����u�6�f�3���/�T`xr�a�%O�w`�!��f�|L;��`�:މ[�xGY;�V�3yn�3����m�c�zN�����1稆���%�u�6�f�3`�f ��{�Hb�0"	ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT������9f?d������D!�yk��	vO���S(�2Y�ǫ�����.���p����o��@(}����ZЖ��ٿE;i���`C>?�{�/z�eg�/�b2�M/��J�W�����ɽ�*<eɽ�*<eɽ�*<e�iƅ���9O�d�!1���s�D�׸ǭ��?��z�IYLy����G8(�2Y�ǫ$W.����|Tu������T�O���ʶ��^�ɽ�*<e��Z0B�񇍞S,��m��8�z4�����iuɽ�*<eɽ�*<eɽ�*<eɽ�*<e�:��MC��;i���`C>�M
��iͮ6s��}�X�
�j�3��9O�d�!1���s�D<��M�D����V��g����j�1���,d������L����^|��]`�W�����ɽ�*<eɽ�*<eɽ�*<e[���g�Q(�2Y�ǫ$W.����|�E��Cӽ��}Mxw��Z0B��3���Kj��˩$�ܚ����t)��`�zN�����1稆���%�u�6�f�3`�f ��{o�Wq�AGɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT������9f?d������&��MS?�)hh�J�.�~��f�|L;��`�:މ[�xGY;�q����d�m`�| ����&�<��f�|L�kC�����o�2��vc �?Y*ɽ�*<eɽ�*<eɽ�*<eɽ�*<e|�'B����u�6�f�3���/�T�A�c���렗k"f+��f�|L;��`�:މ[�xGY;���e�8��������d�zN�����1稆���%�u�6�f�3�Sd�~�fT ��w���7R��ɽ�*<eɽ�*<eɽ�*<e�VJUT������9f?d������$���W 5�m�3'k:�����G8(�2Y�ǫ$W.����|�o�K��o��rK-�'��<��q��M�"���tI�tj�1���,d������Z�?�v&i5%�u�){K۳�EwW�ɽ�*<eɽ�*<eɽ�*<e[���g�Q(�2Y�ǫ$W.����|ar�A�D��^ţ�U�X�
�j�3����N�B�8����竁�F�k	�{d��T��zN�����1稆���%�u�6�f�3�Sd�~�fT ��w���b:n\��ɽ�*<eɽ�*<eɽ�*<e�VJUT������9f?d������aa24얭�@�W�S5�8x�XY��Z0B�񇍞S,��m)��m�.8��l�Ʒ2�v�ɽ�*<e�@����d������Z�?�v&i5Pn���&���!�(I켚<dz�Uiɽ�*<eɽ�*<e[���g�Q(�2Y�ǫ$W.����|ar�A�D��3��|��V8��+ Z5��)ϋ��pᓖC�`E���փ<x@y�07Q���:��e
���4�Qp?��y�ճ���W7P�%(�2Y�ǫ$W.����|�TErǃ+����%֎�5p���ɽ�*<eɽ�*<eɽ�*<e�M,J���ܕpᓖC�6r�?x��}x���Q�˃�6��Rb8�>��z�(�2Y�ǫ$W.����|�o�K��o�E���@��V8��+ Zm`�| �ɽ�*<e��f�|L�kC����m�@�-�F�]��?�`C���z#U�9�ɽ�*<eɽ�*<eɽ�*<e|�'B����u�6�f�3�Sd�~�fTP�d����91��?��!�"
��u�u�6�f�3��ʾ��B`�M�5�쒈��eҥŖqW|9��\ʕpᓖC�`E���փ<�~v3��`@T�;�/ɽ�*<eɽ�*<eɽ�*<e,4���?w��Z0B�񇍞S,��mZm��B��x��kNL�O)ɠo>f��f�|L�kC����pyM��]�|͈��T�<����ZЖ��ٿE;i���`C>?�{�/z���"o��D��Q(�>·�ۃRIɽ�*<eɽ�*<eɽ�*<e�iƅ�����N�B��� @_u}�z�`u�t�,��/;i���`C>?�{�/z���"o��D/��	���Ʒ2�v�ɽ�*<e�@����d������aa24�2G7���"�#F��8��5p���ɽ�*<eɽ�*<e[���g�Q(�2Y�ǫ$W.����|�o�K��o�<�3�N��!�(I�8�>��z�(�2Y�ǫ$W.����|_�_�>_PK"�#F��8S�B���@%����ZЖ��ٿE;i���`C>?�{�/z���"o��D�Z�9�V8��+ Z�W�����ɽ�*<eɽ�*<e�iƅ�����N�B�8���繬d��d��V��P ��Ju9�����Z0B�񇍞S,��m� ��`Rz�6vZ�%�MS�B���@%����Z �jv�5�=�1�ϱ�4��U���5��;#tMɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�1��~!�E�+=�"��~-y75��)ϋ��pᓖC��"��Ѕ�`v�ZP��3_y�|��K[+��1�ϱ������P�۳�EwW�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�1��~!�E�+=�"�����7X�
�j�3����N�BC<ɓ�|*X�i��g��Z�������0{�In<ˋ�DM4Wj̼��Aв�2Gɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��Z0B�񇍞S,��m��eo6����ɒ(�{���	���8���xۄ��\��t\���OxO���<�e�/n<ˋ�DM2�����j�m���[̹ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w�Q�'Ws�t���_��pf��K�`5��)ϋ��pᓖC��"��Ѕ��K�`m`�| �ɽ�*<e�H'b6]�d;+$�.�����d<�8��ЎK�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��~sj@��k����W�Mbg(�!�̸B������;��;i���`C>�M
��iͮf��}J!W-V8��+ Zm`�| �ɽ�*<e�H'b6]�d;+$�.˃�6��Rb�<dz�Uiɽ�*<eɽ�*<eɽ�*<eɽ�*<e��~sj@��k����WJ\O�Z�V8��+ Z5��)ϋ��pᓖC��"��Ѕ�"vЅ\�p;kwֹ���� hyW|9��\�H���5�v����W���P�6;7}x`һaB�ɽ�*<eɽ�*<eɽ�*<e,4���?w��Z0B���Y��� ��j��˩$fMT�Ҁ��O)ɠo>f�/�ӄi�4�kC����k�)�Z�D�Lw��=�zN�����1稆���%I�b�H�`�f ��{I����!�O1�p<�gɽ�*<eɽ�*<eɽ�*<e�VJUT������9f?�(2�oʐSb�&9�ΘQ�z�N̨ <�t-*�5��)ϋ�H���5�Ah�@�;�o��R���7<���^Z�����Ť2��9�|H���5�v����W�������h����&��ɽ�*<eɽ�*<eɽ�*<e,4���?w��Z0B��2h�L�&�_U���)ݝk,�IM�+�I����p�I�b�H�D��}L�8��݌��?ɕ?kV7�hFo+�SZu�L�@�~�>aV�CF�[�
��S�V�堒�c���
��R'ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�/�ӄi�4�kC����=gx�s8�8<�����/�ӄi�4;��`�:މ[�xGY;����8��,*�0�ia�Y�"Woj�1���,�f�� ��E��6��W��#T�m�2��&�ɽ�*<eɽ�*<eɽ�*<e[���g�Q�
T����$W.����| gl�n�!�/��vJ��,d�?���(2�oʐSb�&9��jVYFM�����>W�_��y�ճ���W7P�%�
T����$W.����|�z ��>ԴW�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M,J����H���5�Ah�@�;�o�z �wB���Z0B���Y��� ��j��˩$fMT�Ҁ��m`�| �ɽ�*<e�/�ӄi�4�kC����J��!㣝˻�%e�܉�z�iU�}ɽ�*<eɽ�*<eɽ�*<e|�'B���I�b�H�D��}L�8��݌��?/���?��0�ۧ��5���Z0B��2h�L�&�_,��j��z�IYLy�͵�R}�&ꬶ�RxP�Z�W��
��S�V�堒�c�3�R�3�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�/�ӄi�4�kC�������f�άe[;Zl�fI�b�H�D��}L�8��݌��?;L�?�j7ߔ��� hyW|9��\�H���5�v����W�!&���S+۳�EwW�ɽ�*<eɽ�*<eɽ�*<e,4���?w��Z0B��2h�L�&�_Q�Y�<B�$DX�
�j�3��R~�qB�!1���s�D�|�u�$2���;=6
��y�ճ���W7P�%�
T����$W.����|̃��h�&,m�2��&�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M,J����H���5�Ah�@�;�o�m�[���,d�?���(2�oʐSb�&9��f���ڳ�x�G#�S�t	�g!���j�1���,�f�� ��E��6�J�EL�cm��h�n�gɽ�*<eɽ�*<eɽ�*<e[���g�Q�
T����$W.����|��`��)�:/6�W���,d�?���(2�oʐSb�&9�� kdt]��8���T�JX[��y�ճ���W7P�%�
T����$W.����|�TErǃ++��c��W�����ɽ�*<eɽ�*<eɽ�*<e�M,J����H���5�6r�?x��}x���Q�0�ۧ��5���Z0B��2h�L�&�_Zm��B�R&�[��%q�5�쒈��eҥŖqW|9��\�H���5�ݥ D���z}x���Q���6�Geɽ�*<eɽ�*<eɽ�*<e,4���?w��Z0B��2h�L�&�_)��m�SD+�?M�2D�5�O�I�b�H�Sd�~�fTP�d����8�ꜟ�A��y�ճ���W7P�%�
T����$W.����|�TErǃ+�\�r+�=��W�����ɽ�*<eɽ�*<eɽ�*<e�M,J����H���5�`E���փ<x@y�07Qd!p*�~�X�
�j�3�
��S�V��� @_u}ÙEǛ'�ۄ��\��tZ�����Ť2��9�|H���5�ݥ D���z}x���Q������d<�8��ЎK�ɽ�*<eɽ�*<e,4���?w��Z0B��2h�L�&�_)��m��R�a�G��̸B������;��e���I?�{�/z���"o��D(��Gt�em�B���&��r>�ɽ�*<e��Z0B��2h�L�&�_Ш6�E���f�M�
V8��+ Z�W�����ɽ�*<eɽ�*<e�:��MC��e���I�M
��iͮ���P�V?8����		%Ju9�����Z0B��2h�L�&�_Zm��B�W$�.:�����<���^Q�D@�ɽ�*<e�@�����f��aa24�2G7���7R��ɽ�*<eɽ�*<eɽ�*<e[���g�Q�
T����$W.����|�o�K��o�/�����E�����G8�
T����$W.����|_�_�>_PK�`v�ZP��3_y�|�Mn�_LHw�e���I?�{�/z���"o��D�2nq�Ř�x`һaB�ɽ�*<eɽ�*<eɽ�*<e�iƅ��
��S�V�8���繬d��d��t�T�,G��,d�?���f��$���W 5��;�Y��##m`�| �ɽ�*<e�/�ӄi�4�kC����m�@�-�F��9�:~����7X��q�ɽ�*<eɽ�*<eɽ�*<e|�'B���I�b�H��ʾ��
���B�F�+ ���/�ӄi�4�kC����m�@�-�F�K�@V�sۄ��\��tZ�����Ť2��9�|H���5�`E���փ<�~v3�����'����V8��+ Z�W�����ɽ�*<e,4���?w��Z0B��2h�L�&�_Zm��B��x��kNL������d<�Ju9�����Z0B��2h�L�&�_� ��`Rzǅ؊��SV8��+ Zm`�| �ɽ�*<e�/�ӄi�4�kC����m�@�-�F��I�|�ЮH���<���^�� �R��;ɽ�*<eɽ�*<e|�'B���I�b�H�Sd�~�fTP�d����tseQ,�ٰ���˫�X�
�j�3�
��S�V��� @_u}�r�=_V8��+ Zm`�| �ɽ�*<e�H'b6]{��S�~�!f�� �fɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��~sj@��7f:�El��P�ti+8�̣*���e���I�M
��iͮ9n��5�m`�| ��C4�XȓH'b6]{��S�~��6�Geɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��~sj@��7f:�E���>*�2D�5�O�I�b�H�-�{�0Bh�{"���S����Z �jv�5�=�1�ϱ��Z�F���传]�RH�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�iƅ��
��S�VC<ɓ�|*XS5�8x�XY�Q�'Ws�t�d`�O��P�7rV�܃$����5wz��pN�1�ϱ�D�w*b��v:��Ҟ�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�1��~!E�d�C\���g�@P����H���e���I�M
��iͮ�hc�V�*��Pfɽ�*<e�i�o���Z�I�]�4j�s|Oݽ㺢�"��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����">�{���	���[vC��OG5�td'���ֿ74��/�ӄi�4�kC������7�we*�̸B���Q�D@�ɽ�*<e�i�o���Z�I�]�4���v��{8��ЎK�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����">�{���	���i�(nx�����<���^���;��e���I�M
��iͮO0�-x$�nS�B���@%�܃$���)`���#�`���$��?�{�/z�eg�/�����8�:�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�iƅ��9gi�g !1���s�D�׸ǭ��?�a3#L����,d�?��*��ř%(D!�yk��c�����y�ճ���W7P�%�s7�}��$W.����|�.k-���!!�u�"J�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M,J�����\�m0a�mVW��c�=j0 �M�M�L>�;>cnn37��m�`���$���M
��iͮ�&�ϔ��5�B�������ZЖ��ٿE�`���$��?�{�/z�E�����vL���5ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�iƅ�r)1�ڹ������Cɕ?kV7� 3�/
B�S�s7�}�������.���p�������t�i���+Ȉ4�mJ�KW�B�	E�7;	��7�8`�f ��{�q�
<~�n�C���2ɽ�*<eɽ�*<eɽ�*<e�VJUT������9f?*��ř%(Bx�Ğ��ɘ�n�e�j���,d�?����du�tu�Sb�&9�ΰ��w�]�\\�����v2_�wW|9��\��\�m0a�v����W��Д�٪,�
E�iU�)ɽ�*<eɽ�*<eɽ�*<e,4���?w��Z0B�����V���I��s�$���b\	y`�5��)ϋ��\�m0a�mVW��c�=����E��ݼW��#T���>�K�Rɽ�*<e��Z0B�����V����K��Ɛα,������ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�:��MC�٩`���$���M
��iͮ��s<%��X�
�j�3�9gi�g !1���s�D�׸ǭ��?y*����iɽ�*<e�@����*��ř%(2� ���_d�Ǹ����z#U�9�ɽ�*<eɽ�*<eɽ�*<e[���g�Q�s7�}�������.���p����y�P����g����!�X�
�j�3r)1�ڹ������C/���?��bb����G�zN�����1稆���%;	��7�8`�f ��{�^�WvQt�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT������9f?*��ř%(9v5���6���k��s7�}�������.���p�������/�W�܃$���)`���#�`���$��?�{�/z�k���CЃ�6�Geɽ�*<eɽ�*<eɽ�*<eɽ�*<e�iƅ�r)1�ڹ������Ci���!�)�2D�5�O�;	��7�8D��}L�8��݌��?i���!�)�z�s]eNN`ɽ�*<e��Z0B�����V���X�(��8
c?�4c
�}�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�:��MC�٩`���$���M
��iͮk���C�5��)ϋ��\�m0a�mVW��c�=j0 �MފNf�TJ1rz5���W|9��\��\�m0a�v����W���D�\å@��7�6ɽ�*<eɽ�*<eɽ�*<e,4���?w��Z0B�����V���������t���˾�[(5��)ϋ��\�m0a�mVW��c�=����E���J�EL�cm&��r>�ɽ�*<e��Z0B�����V���Ш6�E���hƁ�,�z�iU�}ɽ�*<eɽ�*<eɽ�*<e�:��MC�٩`���$���M
��iͮ���P�V?��a��{e�X�
�j�3r)1�ڹ��8����竁�F�k	�`v�ZP��3_y�|�Mn�_LHw۩`���$��?�{�/z����P�V?���Jr8�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�iƅ�r)1�ڹ���� @_u}E%��D�&Ը�x-L
��s7�}��$W.����|�o�K��o�Z�H[�MF�z�s]eNN`ɽ�*<e��Z0B�����V���Ш6�E�.8��l·�ۃRIɽ�*<eɽ�*<eɽ�*<e�:��MC�٩`���$��?�{�/z���"o��D�>��y��!�L?7Ƌ;	��7�8��ʾ�� ��w���P�7rV����ZЖ��ٿE�`���$��?�{�/z����P�V?� �^J�����"��ɽ�*<eɽ�*<eɽ�*<e�iƅ�r)1�ڹ���� @_u}����^EG5�td'���ֿ74���?��B��kC����m�@�-�F�L�v:��!�(I�o� ���&ꬶ�RxP�Z�W�r)1�ڹ�yyֶ�T@��PO�K����<���^�� �R��;ɽ�*<eɽ�*<e����n��r��?��B��kC�����V�j��B5+o=�ٰ���˫�X�
�j�3r)1�ڹ��8����竁�F�k	�"vЅ\�p;kwֹZ�����Ť2��9�|�\�m0a�`E���փ<�~v3��>|
ϒ��޴W�����ɽ�*<eɽ�*<e,4���?w��Z0B�����V���Zm��B��x��kNL�0�ۧ��5���Z0B�����V��ؙ ��`Rz�� b��m`�| ���{c^����?��B��kC����m�@�-�F�^�� ���8�:�ɽ�*<eɽ�*<eɽ�*<e|�'B���;	��7�8�Sd�~�fTP�d���ͼ�l�G��5��)ϋ��\�m0a�6r�?x��C'�K��w���� �ɽ�*<e�@����*��ř%(aa24�2G7���b:n\��ɽ�*<eɽ�*<eɽ�*<e[���g�Q�s7�}��$W.����|_�_�>_PK�.���Ȁ���,d�?��*��ř%(aa24�ףr<$�.K�P�7rV����ZЖ��ٿE�`���$��?�{�/z���"o��D j��c�̸B��ຐ �R��;ɽ�*<eɽ�*<e�iƅ�r)1�ڹ��8���繬d��d��ym��Aٰ���˫�X�
�j�3r)1�ڹ���� @_u}c�XO�_ag�̸B���Q�D@�ɽ�*<e�@����*��ř%(aa24�2G7����"vЅ\�����}g�ɽ�*<eɽ�*<e[���g�Q�s7�}��$W.����|�o�K��o����/*� ��K�am@���H�(�;	��7�8��ʾ�֠/��Z �^���<���^Q�D@�ɽ�*<e�i�o�����0>)�k�X P��>d}ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����">�{���	�����j��l��ʏY�u����?��B��kC����]oN�	�L�<��q��M�ZGǦ��4�h}�����0>)�k���5_m��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����">�{���	��S����Ը�x-L
��s7�}��$W.����|r3s��m`�| �ɽ�*<e�H'b6]�)mh�%����QFb�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e|�'B���;	��7�8�-�{�0B;���7d�^���F�*H�4Y����.�NHm`�| ���Da�rF�H'b6]�)mh�%�݁��!8ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��~sj@��R>W�G�^�9	��͟.O@���?��B��kC����5ٗάŻV��X��xB�Z�������0{�I�q �y�Ȍ���\�m�B����h�n�gɽ�*<eɽ�*<eɽ�*<e,4���?w�Q�'Ws�t�^��5"�#F��8k�kN�$���,d�?��*��ř%(���I."lkG5�td'p;kwֹZ�������0{�I�q �y��+��%ƺ��"��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w�Q�'Ws�t�^��5�"vЅ\����ֿ74���?��B��kC����}PYg��?V8��+ Zm`�| �;�e(<�KB�x�#αh�kC����J��!㣝˰T�+Tnɽ�*<eɽ�*<eɽ�*<eɽ�*<e|�'B���@w�����D��}L�8��݌��?/���?��5��)ϋ� �D�O�h>Ah�@�;�o��P�6;7}z�s]eNN`ɽ�*<e��Z0B��>���+�5;~�)�D?R��9����h�n�gɽ�*<eɽ�*<eɽ�*<e�:��MC��m��3+� �IK�vv��8k�>�x��R���7dj�7Y�I�x�#αh�kC�������K�@w� <�t-*�m`�| �ɽ�*<e�x�#αh�kC�����Έx�3�㗟��<�E�W�����ɽ�*<eɽ�*<eɽ�*<e|�'B���@w��������/�T�>��܎�^�7a0b���Z0B�����T|n�j��˩$��}��OI�BDw��?p��y�ճ���Y7W��*�df!п�$W.����|txG�z��h�CÁ�� ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M,J���� �D�O�h>Ah�@�;�o���
���25��)ϋ� �D�O�h>mVW��c�=3��,�����] �, ����Z~�0�V�am��3+� �?�{�/z�wM�.����*��;LAɽ�*<eɽ�*<eɽ�*<eɽ�*<e�iƅ�C�6�vm������C���g�#wf��h�\m��3+� �IK�vv��8k�>�x�Д�٪,�j�M��gt&ꬶ�RxP�Z�W�C�6�vm��堒�c�}�/͓ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�x�#αh�kC����k�)�Z!�"
��u@w�����D��}L�8��݌��?°�:_��Z�����Ť2��9�| �D�O�h>v����W���P�6;7}��H�8�ɽ�*<eɽ�*<eɽ�*<e,4���?w��Z0B�����T|n�j��˩$fMT�Ҁ����T�O�!�"
��u@w��������/�T�f>;�݃f�Ӗ�F>��y�ճ���W7P�%df!п�$W.����|���p�w��W�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M,J���� �D�O�h>Ah�@�;�o�a7���\��Z0B�����T|n�j��˩$&6��u48m`�| �;�e(<�KB�x�#αh�kC�����z��=��3��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e|�'B���@w��������/�TȮ�^q.J1Ը�x-L
�df!п������.���p�����l�06��1	��S��`&ꬶ�RxP�Z�W�C�6�vm��堒�c��[m3Eo�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�x�#αh�kC����(� ��ڷ4-V�]�+ٯm��3+� �IK�vv��8k�>�x�}IU��	����Zq1Q�em��3+� �?�{�/z��QT�G$aW��)f�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�iƅ�C�6�vm������C�[�eonD�Ƣ2�S�m��3+� �IK�vv��8k�>�x��D�\åǓ�Lb�&ꬶ�RxP�Z�W�C�6�vm�yyֶ�T@�����n����z#U�9�ɽ�*<eɽ�*<eɽ�*<e����n��r�x�#αh�kC�����V�j�Mc(J ��!�"
��u@w������Sd�~�fTP�d�����M`.�m`�| ���{c^���x�#αh�kC����K��H7E������W�����ɽ�*<eɽ�*<eɽ�*<e|�'B���@w�������ʾ�� ��w���-��}%����Z0B��>���+�5Zm��B�'y!~ޓ�m1	��S��`&ꬶ�RxP�Z�W�C�6�vm�yyֶ�T@ÙEǛ'��7X��q�ɽ�*<eɽ�*<eɽ�*<e����n��r�x�#αh�kC����m�@�-�F��qA�KJ���
�,��,df!п�$W.����|ar�A�D���\�r+�=�m`�| �ɽ�*<e�x�#αh�kC����K��H7Z�j"�nm�B����h�n�gɽ�*<eɽ�*<e|�'B���@w�������ʾ�� ��w���"�#F��8k�kN�$���,d�?��(�&��aa24얭�@�W������d<�xg��r��*�zN�����1稆���%@w������Sd�~�fT ��w����"vЅ\�����}g�ɽ�*<eɽ�*<e�VJUT������9f?(�&��$���W 5�~��/��K�am@���H�(�@w������Sd�~�fTP�d�������q�ޤS�B���@%����ZЖ��ٿEm��3+� �?�{�/z���"o��D�$@�՛��z�iU�}ɽ�*<eɽ�*<eɽ�*<e�iƅ�C�6�vm��8���繬d��d�2���mX�
�j�3C�6�vm���� @_u}}!�Lڜ<��q��M�"���tI�tj�1���,(�&��aa24�2G7����S�P'qɽ�*<eɽ�*<eɽ�*<e[���g�Qdf!п�$W.����|�o�K��o�����ﴖ=�n\��{Jm��3+� ��M
��iͮ�5�MP���i��g��Z�����Ť2��9�| �D�O�h>`E���փ<�~v3����U������W�����ɽ�*<eɽ�*<e,4���?w��Z0B��>���+�5� ��`RzǍ�����5��)ϋ� �D�O�h>`E���փ<�v�F�
o��U�����m`�| �ɽ�*<e�x�#αh�kC����m�@�-�F�4�)�*�z�G5�td'����}g�ɽ�*<eɽ�*<e|�'B���@w������Sd�~�fTP�d����{M�y0��bm�B�����H�(�@w�������ʾ�֓��P2��G5�td'p;kwֹZ�����Ť2��9�| �D�O�h>`E���փ<�~v3��G������r��5p���ɽ�*<eɽ�*<e,4���?w��Z0B��>���+�5Zm��B��x��kNL�˃�6��Rb8�>��z�df!п�$W.����|_�_�>_PK�"vЅ\�p;kwֹZ�������0{�I9�5P,���X�Y6����F��X
ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w�Q�'Ws�t]1�׮��[��Ur�JF��,d�?��(�&�������1�v�5�쒈�R���%�^����<�e�/9�5P,�}��&�rS�W�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w�Q�'Ws�t]1�׮��-��}%����Z0B��>���+�5�l8�Բ��� �ɽ�*<e�i�o����6�$?���6a�s��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e[���g�Qdf!п�$W.����|+�<b�g�fq�ٓ @�{.6���:��ʵ�~e�Ʒ2�v�!w���y��h}����6�$?��[���MĞ�>υU�%ߏɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����">�{���	�����<�B�����jX.��,d�?��(�&��.���~�$�6��V^�����Z �jv�5�=<�j!l��~�<�_9ұ�!�(I켚<dz�Uiɽ�*<eɽ�*<eɽ�*<eɽ�*<e�1��~!<W��4f%�L�PlC�V8��+ Z5��)ϋ� �D�O�h>�"��Ѕ"�#F��8S�B���@%����Z �jv�5�=<�j!l�������g$$�K�am@���h�n�gɽ�*<eɽ�*<eɽ�*<eɽ�*<e�1��~!<W��4f%��W���k�kN�$���,d�?��(�&��T����=����<���^Q�D@��g����E[��s��kC����J��!㣝˰T�+Tnɽ�*<eɽ�*<eɽ�*<eɽ�*<e[���g�QT��82�9D��}L�8��݌��?/���?��5��)ϋ���;��Y�D!�yk��c�����y�ճ���W7P�%T��82�9`�f ��{I����!�O1�p<�gɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M,J����Ğ(RСܿ�Sb�&9�ΘQ�z�N̨ <�t-*�5��)ϋ���;��Y�&��MS?�)M�L>�;>c���8�ɽ�*<e�愋d�z�kC�����Έx�3�㗟��<�E�W�����ɽ�*<eɽ�*<eɽ�*<e[���g�QT��82�9���/�T�>��܎�^�7a0b��+T��u0������.���p�������t�i���+Ȉ4�mJ�KW�B�	E�7׷�����0�堒�c���
��R'ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���t�$�V'H�kC����=gx�s8�8<�����c�i�#JIK�vv��8k�>�x���
���2m`�| �� ����o�c�i�#J?�{�/z�wM�.����*��;LAɽ�*<eɽ�*<eɽ�*<eɽ�*<e|�'B���׷�����0�����C���g�#wf��h�\E)�dC��mVW��c�=����E��ݼW��#T���>�K�Rɽ�*<e�+T��u0�$W.����|�z ��>ԴW�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�:��MC��E)�dC��Ah�@�;�o�z �wB�+T��u0������.���p����o��@(}����ZЖ��ٿEE)�dC��v����W���P�6;7}��H�8�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e|�Pd]���hӾ�bj��˩$fMT�Ҁ����T�O�!�"
��u׷�����0�����C/���?��bb����G�zN�����1稆���%׷�����0�堒�c�3�R�3�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���t�$�V'H�kC�������f�άe[;Zl�f�Ǐ���J!1���s�D<��M�D����V��g����E[��s��kC�����z��=��3��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e[���g�QT��82�9���/�TȮ�^q.J1Ը�x-L
�T��82�9D��}L�8��݌��?i���!�)�z�s]eNN`ɽ�*<e�+T��u0�$W.����|̃��h�&,m�2��&�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�:��MC��E)�dC��Ah�@�;�o�m�[��w��nR>�;��`�:މ[�xGY;�q����d�m`�| ����&�<�c�i�#J?�{�/z��QT�G$aW��)f�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e|�'B���׷�����0�����C�[�eonD�Ƣ2�S�E)�dC��mVW��c�=����E���J�EL�cm&��r>�ɽ�*<e�+T��u0�$W.����|�TErǃ++��c��W�����ɽ�*<eɽ�*<eɽ�*<e�:��MC��E)�dC��6r�?x��}x���Q�0�ۧ��5��+T��u0�$W.����|�o�K��o��rK-�'��<��q��M�"���tI�tE[��s��kC����K��H7E������W�����ɽ�*<eɽ�*<eɽ�*<e[���g�QT��82�9��ʾ�� ��w���-��}%���+T��u0�$W.����|�o�K��o�Z�H[�MF�z�s]eNN`ɽ�*<e�+T��u0�$W.����|�TErǃ+�\�r+�=��W�����ɽ�*<eɽ�*<eɽ�*<e�:��MC��E)�dC��`E���փ<x@y�07Qd!p*�~�,A�X�>�a���g�_)��m�.8��l�Ʒ2�v�ɽ�*<e�愋d�z�kC����K��H7Z�j"�nm�B����h�n�gɽ�*<eɽ�*<e[���g�QT��82�9��ʾ�� ��w���"�#F��8k�kN�$��w��nR>��kC����m�@�-�F�L�v:��!�(I�o� ���&ꬶ�RqZKǅ�u'a���g�_Ш6�E���f�M�
V8��+ Z�W�����ɽ�*<eɽ�*<e����n��r�c�i�#J�M
��iͮ���P�V?8����		%Ju9���+T��u0�$W.����|�o�K��o�E���@��V8��+ Zm`�| �ɽ�*<e�c�i�#J?�{�/z���"o��D�$@�՛��z�iU�}ɽ�*<eɽ�*<eɽ�*<e|�'B���׷�����0�8���繬d��d�2���m,A�X�>�a���g�_� ��`Rz�� b��m`�| ���{c^�ܘc�i�#J?�{�/z���"o��D�2nq�Ř�x`һaB�ɽ�*<eɽ�*<eɽ�*<e|�'B���׷�����0�8���繬d��d��t�T�,G�w��nR>��kC����pyM��]�|͈��T�<����ZЖ��ٿEE)�dC��`E���փ<�~v3����U������W�����ɽ�*<eɽ�*<eɽ�*<e|�Pd]��a���g�_� ��`RzǍ�����5��)ϋ���;��Y�aa24�ףr<$�.K�P�7rV����ZЖ��ٿEE)�dC��`E���փ<�~v3�����'����V8��+ Z�W�����ɽ�*<eɽ�*<e|�Pd]��a���g�_Zm��B��x��kNL������d<�Ju9���+T��u0�$W.����|_�_�>_PK"�#F��8S�B���@%����ZЖ��ٿEE)�dC��`E���փ<�~v3��G������r��5p���ɽ�*<eɽ�*<eɽ�*<e|�Pd]��a���g�_Zm��B��x��kNL�˃�6��Rb8�>��z�T��82�9��ʾ�֠/��Z �^���<���^Q�D@�ɽ�*<e�i�o���Vnl�@�2�X P��>d}ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����">�{���	��"+[<f�綢ʏY�u���c�i�#J�M
��iͮ9n��5�m`�| ��C4�XȓH'b6]2V���r���6�Geɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��~sj@�#���v���>*�2D�5�O�׷�����0C<ɓ�|*X�i��g��Z�������0{�In!B�dYo4Wj̼��Aв�2Gɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w�+T��u0�$W.����|+�<b�g�fq�ٓ @��#���v:��ʵ�~e�Ʒ2�v�!w���y��h}���Vnl�@�2�[���MĞ�>υU�%ߏɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����">�{���	�����A�Ȅ��jX.�w��nR>��kC����5ٗάŻV��X��xB�Z�������0{�In!B�dYoȌ���\�m�B����h�n�gɽ�*<eɽ�*<eɽ�*<e,4���?w�Q�'Ws�t]a"L���"�#F��8k�kN�$��w��nR>��kC������7�we*�̸B���Q�D@�ɽ�*<e�i�o���Vnl�@�2����v��{8��ЎK�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����">�{���	��a�Z٫����<���^���;��E)�dC���"��Ѕ�"vЅ\�p;kwֹZ������>[��H����G:fGv�{�
;�N�9n��5��W�����ɽ�*<eɽ�*<eɽ�*<e,4���?w���J���:eLE7C<ɓ�|*X0�ۧ��5�	N���^5�}!�Lڜ<��q��M�ZGǦ��4��'�Բ>����q|����7#ub�S�P'qɽ�*<eɽ�*<eɽ�*<eɽ�*<e⃦�q��ڭWH���.a_�A]�l8�Բ�5�8o�-C�f�p�Fv͈��T�<����Z}�����;��F�t�e�&�W�Lƍ3c�3��2·�ۃRIɽ�*<eɽ�*<eɽ�*<eɽ�*<e\<ÌNA�A�1�a��WF�+ ��\���ֻ'��\yJ�	]�� ���ۄ��\��tZ������>[��H����G:fGv�{�
;�N�f��}J!W-V8��+ Z�W�����ɽ�*<eɽ�*<e,4���?w���J���:eLE7C<ɓ�|*X�����d<�Ju9���	N���^5�c�XO�_ag�̸B���Q�D@�ɽ�*<e�� �3Y�S���q|����7#ub�"vЅ\�����}g�ɽ�*<eɽ�*<eɽ�*<e⃦�q��ڭWH���.a_�A]b�l5Q�^�K�am@��� Qoϱm[����v�"vЅ\�p;kwֹZ�����Ť2��9�|2���K,JP�>��7R��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wdFK����f0%ڡV}S�eb����~���}����`�n\#�5�쒈�R���%�^�W|9��\�2���K,JP�>���S�P'qɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wdFK����f0%ڡ�	�D�3%�5�8o�-�|j������k_��=����� �ɽ�*<e��D�MAd ݰm�H�#ڴ-P��7X��q�ɽ�*<eɽ�*<eɽ�*<eɽ�*<erL۪w�Ib}����jk�7�i�F�+ ����7�1��kC�������E-Z�@�Ʒ2�v�ɽ�*<e��D�MAd ݰm�H����v�G5�td'����}g�ɽ�*<eɽ�*<eɽ�*<e[���g�Q����o=$W.����|�e����Ӥm�B���� Qoϱ숨z�<Kc�XO�_ag�̸B���Q�D@�ɽ�*<e��D�MAd ݰm�H+[�&�����<���^�� �R��;ɽ�*<eɽ�*<eɽ�*<e[���g�Q����o=$W.����|cǶcպ��ٰ���˫�9�E虯ء��(���6vZ�%�MS�B���@%����Z��0�)$��|j�����d��ٰ#s�z�iU�}ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e\<ÌNA�'������l>j�m�A����~� e>oGn@al���ɡ�h��b���cTk:�Р˵}�������J�?^�۳�EwW�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<ef��I�����P4�������7A����~� e>oGn@a͈��T�<����Z��0�)$��|j�����.����T�3·�ۃRIɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e\T��}=l[ e>oGn@a�ѥ���ۆ9�E虯�'������M'6/�`��y�ճ��0��hPz8}����"��'L���:��Ҟ�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<ef��I�����P4�����g�@P���}��a�@]�,��pB9Hl�+s���X��xB�Z������&ֵ�0,���a���z��L�PlC�V8��+ Z�W�����ɽ�*<eɽ�*<eɽ�*<e,4���?w��_�'w�R�U�(�N�����d<�Ju9����|P�!�w/ɑ#�����d<�xg��r��*�zN�����(�yi���d;��z�*�+��%ƺ��"��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT��ȏ� P��)?�um��3�	�"vЅ\����ֿ74��E��!�R�wLq?`���<���^Q�D@�ɽ�*<e���'fLSx=��/���K���$5��;#tMɽ�*<eɽ�*<eɽ�*<eɽ�*<e[���g�Q�F{N.J�M
��iͮv�7�w��)�D1��E�)�G��I'�09k� ���ʶ��^��8�
���y|�	R��-L�kC������ޔ��	3x`һaB�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�:��MC��-KB�i��ʾ�֕	�UJو�L�S�ӑ�M�*�%�͈��T�<����ZЖ��ٿE-KB�i�Sd�~�fT����[H\ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e\<ÌNA��¥�c!|�������5��)ϋ�!��QE��j�"c#[tL���ǅҀzN�����1稆���%ҫ�0�7�JP�>��"�#F��8��5p���ɽ�*<eɽ�*<eɽ�*<e�VJUT���e��qb��bSx=��/�J�zܣsT�!�(I��kr���}����7�b��9��G5�td'p;kwֹZ�����Ť2��9�|!��QE����~��!˃�6��Rb�<dz�Uiɽ�*<eɽ�*<eɽ�*<e,4���?w|�	R��-L�kC�����g���pɺV8��+ Z�)�D1��E�)�G��I������^���4�Qp?��y�ճ��vS+ё@}���麲����h��5��;#tMɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<ef��I��鶕)�G��I��~-y7��F9R ���⧼��-�`�n\#�5�쒈�R���%�^����;&�S��SwC˖�A��Vd?o9�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��_�'w�a�eu�^��O)ɠo>f�E��!���e�mꪒr/�0!�$���y�ճ��vS+ё@}����E~���;�_传]�RH�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e���>�(�J�⧼��-�jk�7�i�F�+ ��P���T�Ø(<l�yۄ��\��t\���OxO���;&�S��SwC˖�A���g�@P�M�tb�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��_�'w�a�eu�^��,�o��vA����~��k�P˥��8&ue+�T�!���zN�����(�yi��������y*Ȍ���\�m�B����h�n�gɽ�*<eɽ�*<eɽ�*<e�VJUT��ȏ� P��)?�0�]`~WF"�#F��8k�kN�$ߙ��V�k~�/�Ѭ�c�XO�_ag�̸B���Q�D@�ɽ�*<e���q�Cc�A�`P��"vЅ\�����}g�ɽ�*<eɽ�*<eɽ�*<eɽ�*<erL۪w�Ib}������ȅ�����K�am@� 됰A�k��02v6cD��P�À˃�6��Rbo� ���&ꬶ�RQ�1	�|�-H嵰. ��~��!�!f�� �fɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rIή�%`��kC�����47��W�/t �vwڤBRW/:j��͵�R}��_#��ц2�م|���-H嵰. ��~��!��6�Geɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rIή�%`��kC����t%����|����蛲�@Pek�#0�n �u�HYz�s]eNN`ɽ�*<edFK��Z
�i(�?;�Y�<4~传]�RH�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e1�9 j�*�wڤBRW��6�Q����
�,��,�����x�$W.����|��q�.��9�HF���,ɽ�*<edFK��Z
�i(�?�6S�k�=�!�(I켚<dz�Uiɽ�*<eɽ�*<eɽ�*<e�:��MC��
j����M
��iͮw荦xy�cV8��+ Z�)�D1��E�T�g�MlZp
T�m�B���&��r>�ɽ�*<edFK��Z
�i(�?*?/�=Ȕ�K�am@���h�n�gɽ�*<eɽ�*<eɽ�*<e�:��MC��
j����M
��iͮ��^��Pk�kN�$�L�S�ӑv��g�fDU|M��t+cxg��r��*�zN�����(�yi����M�L�+ҧ�X�Y6����F��X
ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT��ȏ� P��)?'�'�N��q[��Ur�JF���V�k~љ.�;Xb}!�Lڜ<��q��M�ZGǦ��4y�q��^�� ���ƙ�S�P'qɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<erL۪w�Ib}�����N�lܬt�` y氠H����i�~R=�E6�{d��T��zN�����(�yi����M�L�+�4Wj̼��Aв�2Gɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���` �z�U; љ.�;Xb�z�`u�tR?��}�(wڤBRW:��ʵ�~e�Ʒ2�v�!w���y�y�q��^�� ���ƙ��K�`�W�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<erL۪w�Ib}����wl�UoSg�FA��ʗ�|P����MY���u F�yAD*2�&I&ꬶ�R��S����:�pb�j�s|Oݽ㺢�"��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rP���T"t5ů6�	G5�td'���ֿ74��E��!��p�;��XH�؊��SV8��+ Zm`�| �ɽ�*<eP���TtWu�h����<���^�� �R��;ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�"�5ͻ� �@Pek�#0�+��%�ٰ���˫�A����~��R��+��7�D����K�am@�&��r>�ɽ�*<e��Z0B��)�xoĪ���K���$5��;#tMɽ�*<eɽ�*<eɽ�*<eɽ�*<e�:��MC��8�|q{+��M
��iͮv�7�w��)�D1��Em�Y�*��'�09k� ���ʶ��^��8�
���y��Z0B��)�xoĪ�:�W�Ӡ�۳�EwW�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�:��MC��8�|q{+��M
��iͮն��@�fǆ9�E虯ظ�7)�o�+r/�0!�$���y�ճ���W7P�%7��ɇ�F�$W.����|ZO��>t �Aв�2Gɽ�*<eɽ�*<eɽ�*<eɽ�*<ef��I���m�Y�*���I>/�4	�!�L?7Ƌ���H��6��ʾ�����ɃH���y�ճ���W7P�%7��ɇ�F�$W.����|O\�;���m�B����h�n�gɽ�*<eɽ�*<eɽ�*<e�M,J���܇z��X3�
#�k�"�#F��8k�kN�$�L�S�ӑB[�Xs����s��<��G���4�Qp?��y�ճ���W7P�%7��ɇ�F�$W.����||P����J����"��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M,J���܇z��X3�
#�k��"vЅ\����ֿ74�P���TϺ�w���˃�6��Rbo� ���&ꬶ�R��S���l����@�X P��>d}ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rP���T�N�?//�ˢʏY�u���E��!�	j���/Ӹ� b��m`�| ��C4�X�P���T�6�c���,����8�:�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�"�5ͻ� B��Jѻ!�}��&�rS��F9R ���⧼��-��D����A�1	��S��`&ꬶ�R��S���l����@��6a�s��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�E��!�	j���/Ӹ�������)�D1��Em�Y�*�����.�NHm`�| ���Da�rFP���T�H���%j2>��{���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�"�5ͻ� B��Jѻ!�2�����j��y��5}�t�2M�v��g�fDU��BSҧ��H�q/�ɽ�*<e��_�'w���CVD�����d<�8��ЎK�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e1�9 j�*����I�Mbg(�!�̸B�����?-h�j���i�~R�'���5�"�#F��8S�B���@%����Z��0�)$����I��*�jCe�V8��+ Z�W�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<e\<ÌNA� ��P093���v��{Ju9����|P�hsrTq�m������^���4�Qp?��y�ճ���W7P�%RIꐦO�j$W.����|���t������F��X
ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M,J���܁����=�
#�k�[��Ur�JFL�S�ӑ��aE��l���ɡ�h��b���c�)��ן0RIꐦO�j$W.����|uNK�[��ѴW�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M,J���܁����=�
#�k�-��}%����_�'w�w�tF�z���{d��T��zN�����1稆���%�I�\�m�ʹSd�~�fT����[H\ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT��ȏ� P��)?��aE�ũѥ����X�
�j�3^��,Fwpj�"c#[tL���ǅҀzN�����1稆���%�I�\�m�ʹSd�~�fTދF��ݕ���"��ɽ�*<eɽ�*<eɽ�*<e�VJUT������9f?���Lt�c��-��,�ЌG5�td'���ֿ74�P���T�u��:KP�����d<�xg��r��*�zN�����1稆���%�I�\�m�ʹSd�~�fT��9��I�8��ЎK�ɽ�*<eɽ�*<eɽ�*<e�VJUT������9f?���Lt�cߓ�r�\�����<���^��z�v4��B9X�N����7�D����K�am@�&��r>�ɽ�*<e��_�'wڢ�O0�|�!f�� �fɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e1�9 j�*�B9X�N���l��P�ti+�Z��e"����i�~R��`X��`v�ZP��3_y�|��;L���B9X�N����0���Ѓ�x`һaB�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e\<ÌNA���斔�3�&0�w�ڙ��V�k~y��8}v��n �u�HYz�s]eNN`ɽ�*<e��_�'wڢ�O0�|���QFb�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��0'��n���i�~R��`X��.���Ȁ�L�S�ӑ�S���y��P�7rV�܃$���v@-as�3�B9X�N���i�.�!/�pK	��Sɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e\<ÌNA���斔�3�[���MĞ���r1w�6���02v6cϺ�w��¾ƚ�읻�y�ճ��vS+ё@}���麃�F`Z��!�(I켚<dz�Uiɽ�*<eɽ�*<eɽ�*<eɽ�*<ef��I����B_����L�PlC�V8��+ Z��F9R ���⧼��-�zD��IG5�td'p;kwֹZ������&ֵ�0,���_S��`lH��W�����5p���ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��_�'w�m��L�Ӛ�˃�6��Rb�kr���t�2M�B[�Xs���|M��t+cxg��r��*�zN�����1稆���%��+ v���Sd�~�fTɿHd���ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT������9f?��;�T�k�}s�ʏY�u��P���T\=����bb����Gk�w*o��a+O�����+ v���Sd�~�fT��u"+-�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT������9f?��;�T�zÍ�=㓅+�{_R��}�����������1	��S��`&ꬶ�RxP�Z�W�Ɖ�D��0L��~��!���QFb�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rP���T\=����S5�8x�XY��Z0B��n�Rd%��/���M�:~�9�[�P&ꬶ�RxP�Z�W�Ɖ�D��0L��~��!�����d<�8��ЎK�ɽ�*<eɽ�*<eɽ�*<e����n��r;K�Raz�kC�����LJ����]�̸B�����z�v4����4�P�3�|	�!�(I�o� ���&ꬶ�RxP�Z�W�Ɖ�D��0L��~��!˃�6��Rb�<dz�Uiɽ�*<eɽ�*<eɽ�*<e����n��r;K�Raz�kC�����g���pɺV8��+ Z�)�D1��E<�a�a�������^���4�Qp?��y�ճ��vS+ё@}�������b6�H5��;#tMɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<ef��I���<�a�a맾�~-y7��F9R ���⧼��-�?KErB��'�5�쒈�R���%�^����;&�S����QkK��Vd?o9�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��_�'w��?*�ڡ��O)ɠo>f�E��!��8�טCv�r/�0!�$���y�ճ��vS+ё@}����cA���wF传]�RH�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e���>�(�J�⧼��-�4�H�LFF�+ ��P���T��2b>[m�ۄ��\��t\���OxO���;&�S����QkK���g�@P�M�tb�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��_�'w��?*�ڡ��,�o��vA����~�����>>���8&ue+�T�!���zN�����(�yi����ߕ�)���Ȍ���\�m�B����h�n�gɽ�*<eɽ�*<eɽ�*<e�VJUT��ȏ� P��)?C�ypVq�"�#F��8k�kN�$ߙ��V�k~�%�,K/�>c�XO�_ag�̸B���Q�D@�ɽ�*<e���q�Cs��ĵ��&�"vЅ\�����}g�ɽ�*<eɽ�*<eɽ�*<eɽ�*<erL۪w�Ib}�����#w}tܺ�K�am@� 됰A�k��02v6c�u��:KP˃�6��Rbo� ���&ꬶ�RxP�Z�W�q>��Z�.���~��!�!f�� �fɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r��3����kC�����47��W�/t �v0 A��!M/:j��͵�R}��_#��ц2aV�CF�[q>��Z�.���~��!��6�Geɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r��3����kC����t%����|����蛲w	z9��蹤n �u�HYz�s]eNN`ɽ�*<e��Z0B��N'�����;�Y�<4~传]�RH�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e1�9 j�*�0 A��!M��6�Q����
�,��,�ϝO�}�$W.����|��q�.��9�HF���,ɽ�*<e��Z0B��N'������6S�k�=�!�(I켚<dz�Uiɽ�*<eɽ�*<eɽ�*<e�:��MC��|m9T�g�R�M
��iͮw荦xy�cV8��+ Z�)�D1��E#vw8���MlZp
T�m�B���&��r>�ɽ�*<e��Z0B��N'�����*?/�=Ȕ�K�am@���h�n�gɽ�*<eɽ�*<eɽ�*<e�:��MC��|m9T�g�R�M
��iͮ��^��Pk�kN�$�L�S�ӑ�fC&u�|M��t+cxg��r��*�zN�����(�yi����c���b��X�Y6����F��X
ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT��ȏ� P��)?���_��pf[��Ur�JF���V�k~��C�jli�}!�Lڜ<��q��M�ZGǦ��4y�q��^����ܠ�X��S�P'qɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<erL۪w�Ib}����'�H�����` y氠H����i�~R��񤿶`)�{d��T��zN�����(�yi����c���b4Wj̼��Aв�2Gɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���` �z�U; ��C�jli��z�`u�tR?��}�(0 A��!M:��ʵ�~e�Ʒ2�v�!w���y�y�q��^����ܠ�X���K�`�W�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<erL۪w�Ib}����U������g�FA��ʗ�|Pӡ�I;P��E�u F�yAD*2�&I&ꬶ�R��S����D����vHj�s|Oݽ㺢�"��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rP���T�!�,�ǁG5�td'���ֿ74��E��!��h��S�Յ؊��SV8��+ Zm`�| �ɽ�*<eP���T��!T �����<���^�� �R��;ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�"�5ͻ� w	z9����+��%�ٰ���˫�A����~�|�>��~�7�D����K�am@�&��r>�ɽ�*<e��Z0B�񇍞S,��m���K���$5��;#tMɽ�*<eɽ�*<eɽ�*<eɽ�*<e�:��MC��;i���`C>�M
��iͮv�7�w��)�D1��E��������'�09k� ���ʶ��^��8�
���y��Z0B�񇍞S,��m�:�W�Ӡ�۳�EwW�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�:��MC��;i���`C>�M
��iͮն��@�fǆ9�E虯�,E�}PO��r/�0!�$���y�ճ���W7P�%(�2Y�ǫ$W.����|ZO��>t �Aв�2Gɽ�*<eɽ�*<eɽ�*<eɽ�*<ef��I��鶤��������I>/�4	�!�L?7Ƌ�u�6�f�3��ʾ�����ɃH���y�ճ���W7P�%(�2Y�ǫ$W.����|O\�;���m�B����h�n�gɽ�*<eɽ�*<eɽ�*<e�M,J���ܕpᓖC�
#�k�"�#F��8k�kN�$�L�S�ӑbO�1��	��s��<��G���4�Qp?��y�ճ���W7P�%(�2Y�ǫ$W.����||P����J����"��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M,J���ܕpᓖC�
#�k��"vЅ\����ֿ74�P���T��9�x˃�6��Rbo� ���&ꬶ�R��S�������f:�X P��>d}ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rP���T�����9ǢʏY�u���E��!�<���`<T� b��m`�| ��C4�X�P���T�AY��������8�:�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�"�5ͻ� 1bF��E߈}��&�rS��F9R ���⧼��-�CvG�j8O1	��S��`&ꬶ�R��S�������f:��6a�s��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�E��!�<���`<T�������)�D1��E�����������.�NHm`�| ���Da�rFP���T�/V ���/2>��{���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�"�5ͻ� 1bF��E߈2�����j��y��5}�t�2M��fC&u���BSҧ��H�q/�ɽ�*<e��_�'w�{��S�~�����d<�8��ЎK�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e1�9 j�*�|���%
�Mbg(�!�̸B�����?-h�j���i�~R��) �"�#F��8S�B���@%����Z��0�)$�|���%
��*�jCe�V8��+ Z�W�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<e\<ÌNA��Ҙp�f�����v��{Ju9����|PӫE�+=�"������^���4�Qp?��y�ճ���W7P�%�
T����$W.����|���t������F��X
ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M,J����H���5�
#�k�[��Ur�JFL�S�ӑ J^���l���ɡ�h��b���c�)��ן0�
T����$W.����|uNK�[��ѴW�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M,J����H���5�
#�k�-��}%����_�'w�$`��`W�{d��T��zN�����1稆���%I�b�H�Sd�~�fT����[H\ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT��ȏ� P��)? J^����ѥ����X�
�j�3�
��S�Vj�"c#[tL���ǅҀzN�����1稆���%I�b�H�Sd�~�fTދF��ݕ���"��ɽ�*<eɽ�*<eɽ�*<e�VJUT������9f?�f���-��,�ЌG5�td'���ֿ74�P���T�K��(��à����d<�xg��r��*�zN�����1稆���%I�b�H�Sd�~�fT��9��I�8��ЎK�ɽ�*<eɽ�*<eɽ�*<e�VJUT������9f?�f����r�\�����<���^��z�v4��sKh��dT�7�D����K�am@�&��r>�ɽ�*<e��_�'w��)mh�%��!f�� �fɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e1�9 j�*�sKh��dTl��P�ti+�Z��e"����i�~Rh���h�E�`v�ZP��3_y�|��;L���sKh��dT�0���Ѓ�x`һaB�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e\<ÌNA��)Y[���j&0�w�ڙ��V�k~)T��ׄHT�n �u�HYz�s]eNN`ɽ�*<e��_�'w��)mh�%����QFb�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��0'��n���i�~Rh���h�E�.���Ȁ�L�S�ӑ�^��5�P�7rV�܃$���v@-as�3�sKh��dTi�.�!/�pK	��Sɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e\<ÌNA��)Y[���j[���MĞ���r1w�6���02v6c��9�x�ƚ�읻�y�ճ��vS+ё@}�����I	�FHA��!�(I켚<dz�Uiɽ�*<eɽ�*<eɽ�*<eɽ�*<ef��I��鶳@E�CS��L�PlC�V8��+ Z��F9R ���⧼��-������R�G5�td'p;kwֹZ������&ֵ�0,��oC�K$�����W�����5p���ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��_�'wڲ��;~*�˃�6��Rb�kr���t�2M�bO�1��	�|M��t+cxg��r��*�zN�����1稆���%;	��7�8�Sd�~�fTɿHd���ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT������9f?*��ř%(�k�}s�ʏY�u��P���T?�R�ף�bb����Gk�w*o��a+O���;	��7�8�Sd�~�fT��u"+-�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT������9f?*��ř%(�zÍ�=㓅+�{_R���g�ʿ�Ϲ|�q�u �1	��S��`&ꬶ�RxP�Z�W�r)1�ڹ���~��!���QFb�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rP���T?�R�ף�S5�8x�XY��Z0B�����V����/���M�:~�9�[�P&ꬶ�RxP�Z�W�r)1�ڹ���~��!�����d<�8��ЎK�ɽ�*<eɽ�*<eɽ�*<e����n��r��?��B��kC�����LJ����]�̸B�����z�v4���U��_��P�3�|	�!�(I�o� ���&ꬶ�RxP�Z�W�r)1�ڹ���~��!˃�6��Rb�<dz�Uiɽ�*<eɽ�*<eɽ�*<e����n��r��?��B��kC�����g���pɺV8��+ Z�)�D1��Ei�27�?p�������^���4�Qp?��y�ճ��vS+ё@�g�ʿ�Ϲ��$i8�5��;#tMɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<ef��I���i�27�?p���~-y7��F9R ���⧼��-�Ը��!��5�쒈�R���%�^����;&�S���(ϰ�Y���Vd?o9�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��_�'w�Y/�P`�&�O)ɠo>f�E��!��y�k	o6r/�0!�$���y�ճ��vS+ё@�g�ʿ�Ϲ������R�传]�RH�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e���>�(�J�⧼��-��}Mu?�F�+ ��P���T�K�L�+b�ۄ��\��t\���OxO���;&�S���(ϰ�Y����g�@P�M�tb�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��_�'w�Y/�P`�&�,�o��vA����~�L2�*<*SͰ�8&ue+�T�!���zN�����(�yi���>��@��8�Ȍ���\�m�B����h�n�gɽ�*<eɽ�*<eɽ�*<e�VJUT��ȏ� P��)?]1�׮��"�#F��8k�kN�$ߙ��V�k~�/�����c�XO�_ag�̸B���Q�D@�ɽ�*<e���q�C�� �O��"vЅ\�����}g�ɽ�*<eɽ�*<eɽ�*<eɽ�*<erL۪w�Ib�g�ʿ�ϹDB�hDx3�K�am@� 됰A�k��02v6c�K��(���˃�6��Rbo� ���&ꬶ�RxP�Z�W�C�6�vm���~��!�!f�� �fɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�x�#αh�kC�����47��W�/t �vD�Ɂ�p��/:j��͵�R}��_#��ц2aV�CF�[C�6�vm���~��!��6�Geɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�x�#αh�kC����t%����|����蛲X��0/�Фn �u�HYz�s]eNN`ɽ�*<e��Z0B��>���+�5;�Y�<4~传]�RH�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e1�9 j�*�D�Ɂ�p����6�Q����
�,��,df!п�$W.����|��q�.��9�HF���,ɽ�*<e��Z0B��>���+�5�6S�k�=�!�(I켚<dz�Uiɽ�*<eɽ�*<eɽ�*<e�:��MC��m��3+� ��M
��iͮw荦xy�cV8��+ Z�)�D1��E/i	�ꐔ�MlZp
T�m�B���&��r>�ɽ�*<e��Z0B��>���+�5*?/�=Ȕ�K�am@���h�n�gɽ�*<eɽ�*<eɽ�*<e�:��MC��m��3+� ��M
��iͮ��^��Pk�kN�$�L�S�ӑ�����p�
|M��t+cxg��r��*�zN�����(�yi���������駣X�Y6����F��X
ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT��ȏ� P��)?]a"L���[��Ur�JF���V�k~NvX���_�}!�Lڜ<��q��M�ZGǦ��4y�q��^�ŃQZ1���S�P'qɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<erL۪w�Ib�g�ʿ�Ϲ�&*A��~]` y氠H����i�~R��YjI]�{d��T��zN�����(�yi����������4Wj̼��Aв�2Gɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���` �z�U; NvX���_��z�`u�tR?��}�(D�Ɂ�p��:��ʵ�~e�Ʒ2�v�!w���y�y�q��^�ŃQZ1����K�`�W�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<erL۪w�Ib�g�ʿ�Ϲ���|�zg�FA��ʗ�|P�<W��4f%�u F�yAD*2�&I&ꬶ�R��S������9?�YAj�s|Oݽ㺢�"��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rP���T��9�5yG5�td'���ֿ74��E��!�c�����؊��SV8��+ Zm`�| �ɽ�*<eP���T�s*���|���<���^�� �R��;ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�"�5ͻ� X��0/���+��%�ٰ���˫�A����~��d-0�Ų�7�D����K�am@�&��r>�ɽ�*<e�+T��u0�$W.����|���t������F��X
ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�:��MC��E)�dC��
#�k�[��Ur�JFL�S�ӑ�o2 U�Y�l���ɡ�h��b���c�)��ן0T��82�9�Sd�~�fT��u"+-�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M,J������;��Y��zÍ�=㓅+�{_R���g�ʿ�ϹyZ�͂�1	��S��`&ꬶ�RqZKǅ�u'a���g�_;�Y�<4~传]�RH�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rP���Tx>��e���S5�8x�XY�+T��u0�$W.����|��q�.��9�HF���,ɽ�*<e�+T��u0�$W.����|O\�;���m�B����h�n�gɽ�*<eɽ�*<eɽ�*<e�:��MC��E)�dC��
#�k�"�#F��8k�kN�$�L�S�ӑ�o2 U�Y��s��<��G���4�Qp?��y�ճ���W7P�%T��82�9�Sd�~�fT��9��I�8��ЎK�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�M,J������;��Y���r�\�����<���^��z�v4����e����7�D����K�am@�&��r>�ɽ�*<e��_�'w�8�'	ϛ�i�!f�� �fɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e1�9 j�*���e���l��P�ti+�Z��e"����i�~R~��V�E��`v�ZP��3_y�|��;L�����e����0���Ѓ�x`һaB�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e\<ÌNA�8a����&0�w�ڙ��V�k~p������n �u�HYz�s]eNN`ɽ�*<e��_�'w�8�'	ϛ�i���QFb�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��0'��n���i�~R~��V�E��.���Ȁ�L�S�ӑ��-t邜P�7rV�܃$���v@-as�3���e���i�.�!/�pK	��Sɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e\<ÌNA�8a����[���MĞ���r1w�6���02v6c�s{8�9���ƚ�읻�y�ճ��vS+ё@�g�ʿ�Ϲa�9�5���!�(I켚<dz�Uiɽ�*<eɽ�*<eɽ�*<eɽ�*<ef��I���K����J���L�PlC�V8��+ Z��F9R ��`m�J�d�< �\��G5�td'p;kwֹZ������&ֵ�0,��W-���zӡ�W�����5p���ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��_�'w��D�����&˃�6��Rb�kr���t�2M������p�
|M��t+cxg��r��*�zN�����(�yi���B��$�J�!f�� �fɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT��ȏ� P��)?l��P�ti+������F�t�e�W���ߺ���y����}!�Lڜ<��q��M�ZGǦ��4y�q��^��0���Ѓ�x`һaB�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<erL۪w�Ib�r��z�>1&0�w��|��z8�2���q|���TQF�ڗ_(�S�����{d��T��zN�����(�yi���B��$�J���QFb�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���M�{�Z����q|���TQF�ڗ_(�S�����.���Ȁ�L�S�ӑ:��ʵ�~e�Ʒ2�v�!w���y�y�q��^�i�.�!/�pK	��Sɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<erL۪w�Ib�r��z�>1[���MĞ�μ�4���j��Ehf�+3yH&0�a�N�u F�yAD*2�&I&ꬶ�R��S�������"��!�(I켚<dz�Uiɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�0_�����L�PlC�V8��+ Zi �Dl�<O�G:fGv��Y����#RC��y�؊��SV8��+ Zm`�| �ɽ�*<e�#��w���W�����5p���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�"�5ͻ� �
(��c�˃�6��Rb��3h5�DڭWH��3�A�f<��SOC�u��J7�����K�am@�&��r>��8�
���y���J�����XPs�P2�0x����&�P������8�:�ɽ�*<eɽ�*<eɽ�*<eX�T.6���F�t�e�W���ߺ���y����}��&�rS�F����[Gm��g�r/�0!�$���y�ճ��8�1���E�ڭWH��3�A�f<��T�;��.����T�3·�ۃRIɽ�*<eɽ�*<eɽ�*<e!��$и3�[Gm��g�������i �Dl�<O�G:fGv��Y����#.cu,"y�zM'6/�`��y�ճ��
�_�ڭWH��3�A�f<��T�;��i�.�!/�pK	��Sɽ�*<eɽ�*<eɽ�*<e\�@?<���G:fGv��Y����#.cu,"y�z[���MĞ���kg@0���4B�-�u F�yAD*2�&I&ꬶ�R�E�HP8jΗCf�|��$EB<b���L�"�#F��8��5p���ɽ�*<eɽ�*<e����n��r\���ֻ'�[\r�R��&��J!���U��+�r�!�(I�"j��5����=a�^�P�3�|	�!�(I�o� ���&ꬶ�R�E�HP8jΗCf�|��$EB<b���L��"vЅ\�����}g�ɽ�*<eɽ�*<e����n��r\���ֻ'�[\r�R��&��J!�����?Պl�K�am@�F�c�0.-��4B�-������^���4�Qp?��y�ճ��vS+ё@Z���^S��~-y7�W�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e���>�(�J�za[��[�0�ۧ��5����J�����XPs�P'��LE��2��z�bb����Gk�w*o�Ё]-Ԗ���׈{w�J�S�P'qɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���}�B-u����/<�k�?a�G���F�t�e�W���ߺ�)����36�n �u�HYz�s]eNN`ɽ�*<e�ƾYn��d.����T�3·�ۃRIɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eX�T.6���F�t�e�W���ߺ�)����36�z�`u�t���	�9t�t���M'6/�`��y�ճ��0��hPz8Z���^S���g�@P�M�tb�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e���>�(�J�za[��[�,�o��v����pQcΗCf�|��$EB<b��.����$��BSҧ��H�q/�ɽ�*<e�ƾYn��d!`h FH�
�̸B��ຐ �R��;ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��0'��n�t���j�s|Oݽ�ٰ���˫����pQcΗCf�|��$EB<b��.����$�s��<��G���4�Qp?��y�ճ��vS+ё@Z���^S��W�����5p���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e���>�(�J�za[��[�˃�6��Rb��3h5�DڭWH��3�A�f<���p��Ar�J7�����K�am@�&��r>�ɽ�*<e���J�����XPs�P�Ĝ�9�%,�ydb�=��z#U�9�ɽ�*<eɽ�*<eɽ�*<eX�T.6���F�t�e�W���ߺ�)����36��X�Y6�B��焷sm�j��Eh_����ncܖ�	ǯJ��ʶ��^��8�
���y���J�����XPs�P�Ĝ�9�%�����В���8�:�ɽ�*<eɽ�*<eɽ�*<eX�T.6���F�t�e�W���ߺ�)����36}��&�rSi �Dl�<O�G:fGv���=HD����T9O�3Y��y�ճ��8�1���E�ڭWH��3�A�f<㋞�TUn��.����T�3·�ۃRIɽ�*<eɽ�*<eɽ�*<e\�@?<���G:fGv���=HD���(��ʸG�i �Dl�<O�G:fGv��Y����#ј>�^�M'6/�`��y�ճ��
�_�ڭWH��3�A�f<㋞�TUn��i�.�!/�pK	��Sɽ�*<eɽ�*<eɽ�*<e\�@?<���G:fGv��Y����#ј>�^�[���MĞ�μ�4���j��Eh_����nc{"g/R�AD*2�&I&ꬶ�R�E�HP8jΗCf�|��$EB<b eE���A�"�#F��8��5p���ɽ�*<eɽ�*<e����n��r\���ֻ'�[\r�R���?�9⻔��̢���k�!�(I���3h5�DڭWH���.a_�A]�J�zܣsT�!�(I�o� ���&ꬶ�R�E�HP8jΗCf�|��$EB<b eE���A��"vЅ\�����}g�ɽ�*<eɽ�*<e����n��r\���ֻ'�[\r�R���?�9⻔�K�-}�J�K�am@�1�~46΋@�j��Eh_����nccǶcպ�����4�Qp?��y�ճ��:j���+���=a�^��) �)x5��;#tMɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e!��$и3�|��@S��jME���:�F����*/1Fu=S&��ؒh��b���c��Gj�B�����=a�^����@�^�۳�EwW�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e!��$и3�|��@S��x����s��^����0�n	���{d��T��zN������%,!u�r�u^jP��:旿�]��Aв�2Gɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���Օ�^�e�L*S5�8x�XY�7cϢA����<&0~L���ǅҸL�~bq�}�qТ�j�u^jP��:�;������m���[̹ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT��ȅV�)��C�a�jN<��K�`�F����*/1Fu=S�8����c��H�q/�ɽ�*<e�7cϢA�f;��@�!�����d<�8��ЎK�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��S�"��[�#�Vxg��}ɻ�&lc�̸B���R�:�`�<�<��m�ƿy��>��m�B���&��r>�ɽ�*<e�7cϢA�f;��@�!˃�6��Rb�<dz�Uiɽ�*<eɽ�*<eɽ�*<eɽ�*<e��S�"��[�#�Vxg�>5xW�V8��+ Z�F����*/1Fu=S}<��m�xg��r��*�zN������%,!u�r�u^jP��:���R�8
����F��X
ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT��ȅV�)��w��Z�[��Ur�JFj�����e�mꪒ}�1�|�0c��ʶ��^��8�
���y�7cϢA�F��y��6�Geɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��S�"��[�#�Vxg�g��E{j���
��E�	c�W.�ҽ�E��9 1	��S��`&ꬶ�R��<nK&�_�,�\���8����V_ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�H'b6]C���-!����� �$Q��z�X����N$ݯ`��y�׻�y�ճ��`#�F�\���=a�^&�i���:��Ҟ�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e!��$и3�|��@S���8D��t����xE�}�1�ϱ��3)��q�ƚ�읻�y�ճ��:j���+���=a�^
0��Y~�!�(I켚<dz�Uiɽ�*<eɽ�*<eɽ�*<eɽ�*<e!��$и3�|��@S��}�g9�bV8��+ Z�F����/�Ѭ����'�1�!�(I�o� ���&ꬶ�R��<nK&�_�,�\���F�x�N8��ЎK�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r1�"�-�d�y������<���^R�:�`�<�1�ϱ��3)��q˃�6��Rbo� ���&ꬶ�R��<nK&�_�,�\�����W�
�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r1�"�-��k3�8��ʏY�u���H'b6]=�E6&��ؒh��b���c��Gj�B�����=a�^�]���b�۳�EwW�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e!��$и3�|��@S��d� ��Y���^������MY��KlR41uz�s]eNN`ɽ�*<e�7cϢA�u�?[)������QFb�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��S�"���1�ϱ���i�,2ES5�8x�XY�7cϢA�fD1�3�L���ǅҸL�~bq�}�qТ�j�u^jP��:�铫h�m���[̹ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT��ȅV�)��J�m@��K�`�F����љ.�;Xb� O�bë�T�!���zN������%,!u�r�u^jP��:�����2@m�B����h�n�gɽ�*<eɽ�*<eɽ�*<e�VJUT��ȅV�)��J�m@"�#F��8k�kN�$�j������p�;��XHy��>��m�B���&��r>�ɽ�*<e�7cϢA�u�?[)���˃�6��Rb�<dz�Uiɽ�*<eɽ�*<eɽ�*<eɽ�*<e��S�"��[�#�Vxg�V��Y�DPV8��+ Z�F����љ.�;Xb�RC^��K�am@�&��r>�ɽ�*<e�7cϢA���4ŭE�B�!f�� �fɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��S�"��[�#�Vxg��T�7�3�	.�v���T��1�ϱ�Wd���UɆbb����Gk�w*o�=��wY��u^jP��:[��|S��%�W�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT��ȅV�)�VϚ&L��-��}%���Q�'Ws�tv��g�fDU�ӝE+<�u��y�ճ��:j���+���=a�^�OU��Dۀ传]�RH�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e!��$и3��:��*�Ɛ�sg���ɒ(夜��=a�^�ξ���:~�9�[�P9��7�rXS��<�#l�_�,�\����|���I�>υU�%ߏɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r1�"�-2�0��|S���jX.j������	j���/Ӹ�5� 2�9AD*2�&I&ꬶ�R��<nK&�_�,�\��xξ>�f���"��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r1�"�-!>\�����G5�td'���ֿ74ēH'b6]�'���5�8�� �a����4�Qp?��y�ճ��:j���+���=a�^��.;7㳮�K�am@���h�n�gɽ�*<eɽ�*<eɽ�*<eɽ�*<e!��$и3�|��@S��&Py�eH�k�kN�$�j������	j���/Ӹ|Gb��f	>���4�Qp?��y�ճ��:j���+���=a�^$��HP��5��;#tMɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e!��$и3�|��@S��ZF����\�F����y��8}v�©�U>�T@�͵�R}��_#��ц2XS��<�#l�_�,�\��^��e|��9ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r1�"�-,<�~:���#��c���H{���	������.��R�{d��T��zN������%,!u�r�u^jP��:&�Ջ��`
Aв�2Gɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���Օ�^�e��,�⮾�[��p��q�ٓ @���4B�-&�Ջ��`
9�HF���,u�)�P�7cϢA��`�j�Y�i݁��!8ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��S�"��[�#�Vxg���8��Q��͟.O@��H'b6]��`X��8����c��H�q/�ɽ�*<e�7cϢA��`�j�Y�i�����d<�8��ЎK�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��S�"��[�#�Vxg�l}ڞ9mx>�̸B���R�:�`�<�1�ϱ�Ģ��0$�����d<�xg��r��*�zN������%,!u�r�u^jP��:��&qƕ���"��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT��ȅV�)��t;Yi���"vЅ\����ֿ74ēH'b6]��`X�}<��m�xg��r��*�zN������%,!u�r�u^jP��:�'��pD	۵��F��X
ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT��ȅV�)�XqLU:M[��Ur�JFj������8�טCv�}�1�|�0c��ʶ��^��8�
���y�7cϢA�ꗡ��E����6�Geɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��S�"��[�#�Vxg�;NM�4e��
��E�
	}�%I�E��9 1	��S��`&ꬶ�R��<nK&�_�,�\���pE�xt�Qɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�H'b6]w�tF�z��!����� �$Q��z�X����N$���9?Ga���y�ճ��`#�F�\���=a�^J<N���(.:��Ҟ�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e!��$и3�|��@S��5����Վ��xE�}�1�ϱ����,�l�ƚ�읻�y�ճ��:j���+���=a�^_^3���!�(I켚<dz�Uiɽ�*<eɽ�*<eɽ�*<eɽ�*<e!��$и3�|��@S����!@%XrV8��+ Z�F����%�,K/�>���'�1�!�(I�o� ���&ꬶ�R��<nK&�_�,�\���<sEvT8��ЎK�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r1�"�-P��9W�|���<���^R�:�`�<�1�ϱ����,�l˃�6��Rbo� ���&ꬶ�R��<nK&�_�,�\���67�lȿɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r1�"�-`��'��ʏY�u���H'b6]��񤿶`)&��ؒh��b���c��Gj�B�����=a�^t&*���	�۳�EwW�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e!��$и3�|��@S���z�c*���^�����I;P��EKlR41uz�s]eNN`ɽ�*<e�7cϢA�jQ��օ�����QFb�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��S�"���1�ϱ�u)n�	�	�S5�8x�XY�7cϢA�����9��}L���ǅҸL�~bq�}�qТ�j�u^jP��:������;m���[̹ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT��ȅV�)�74P�=ā��K�`�F�����C�jli�� O�bë�T�!���zN������%,!u�r�u^jP��:�zH�8��m�B����h�n�gɽ�*<eɽ�*<eɽ�*<e�VJUT��ȅV�)�74P�=ā"�#F��8k�kN�$�j������h��S��y��>��m�B���&��r>�ɽ�*<e�7cϢA�jQ��օ��˃�6��Rb�<dz�Uiɽ�*<eɽ�*<eɽ�*<eɽ�*<e��S�"��[�#�Vxg����7��w�V8��+ Z�F�����C�jli��RC^��K�am@�&��r>�ɽ�*<e�7cϢA��_P���a��!f�� �fɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��S�"��[�#�Vxg�����c�.�v���T��1�ϱ���pd��cbb����Gk�w*o�=��wY��u^jP��:ԟ|��{��W�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT��ȅV�)���T����-��}%���Q�'Ws�t�fC&u��ӝE+<�u��y�ճ��:j���+���=a�^����B!"传]�RH�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e!��$и3���=�*�ꚯƐ�sg���ɒ(夜��=a�^��]�|w�q:~�9�[�P9��7�rXS��<�#l�_�,�\���� !!>υU�%ߏɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r1�"�-~T�<2���jX.j������<���`<T�5� 2�9AD*2�&I&ꬶ�R��<nK&�_�,�\���>���cº��"��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r1�"�-sb(�ZG5�td'���ֿ74ēH'b6]��) �8�� �a����4�Qp?��y�ճ��:j���+���=a�^�d��X(
�K�am@���h�n�gɽ�*<eɽ�*<eɽ�*<eɽ�*<e!��$и3�|��@S��x`�Yk�kN�$�j������<���`<T|Gb��f	>���4�Qp?��y�ճ��:j���+���=a�^:J��]��5��;#tMɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e!��$и3�|��@S���)�`?i��F����)T��ׄHT©�U>�T@�͵�R}��_#��ц2XS��<�#l�_�,�\���u@��M�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r1�"�-�/�����#��c���H{���	������W'�{d��T��zN������%,!u�r�u^jP��:z#�*C�M1Aв�2Gɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���Օ�^�e�gB���[��p��q�ٓ @���4B�-z#�*C�M19�HF���,u�)�P�7cϢA��)[���/f݁��!8ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��S�"��[�#�Vxg���qje�.0�͟.O@��H'b6]h���h�E�8����c��H�q/�ɽ�*<e�7cϢA��)[���/f�����d<�8��ЎK�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��S�"��[�#�Vxg�Lͼr�!�̸B���R�:�`�<�1�ϱ�w�����������d<�xg��r��*�zN������%,!u�r�u^jP��:�w��������"��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT��ȅV�)�mT����Tv�"vЅ\����ֿ74ēH'b6]h���h�E}<��m�xg��r��*�zN������%,!u�r�u^jP��:��>9S���F��X
ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT��ȅV�)���Ǽ��x[��Ur�JFj������y�k	o6}�1�|�0c��ʶ��^��8�
���y�7cϢA����j�� ��6�Geɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��S�"��[�#�Vxg������mà��
��E���R>W�G��E��9 1	��S��`&ꬶ�R��<nK&�_�,�\������V3�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�H'b6]$`��`W!����� �$Q��z�X����N$݀��X-�����y�ճ��`#�F�\���=a�^�P�����$:��Ҟ�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e!��$и3�|��@S��ٳ:�W�����xE�}�1�ϱ�\�y1Sa�ƚ�읻�y�ճ��:j���+���=a�^Ӿ��h��!�(I켚<dz�Uiɽ�*<eɽ�*<eɽ�*<eɽ�*<e!��$и3�|��@S��]T�� [V8��+ Z�F����/��������'�1�!�(I�o� ���&ꬶ�R��<nK&�_�,�\��t�99�`��8��ЎK�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r1�"�-t߶j\�j���<���^R�:�`�<�1�ϱ�\�y1Sa˃�6��Rbo� ���&ꬶ�R��<nK&�_�,�\��]R�z�.k�W�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r1�"�-����m��0�ۧ��5��Q�'Ws�tʨ��ehz�i� P�m`�| ��C4�X�1�"�-�U���Q��6�Geɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��~sj@��4B�-$$p�X�Ҷ��
��E�{.6����E��9 1	��S��`&ꬶ�R��<nK&�_�,�\���앫�;`p�W�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�H'b6]��YjI]!����� �$Q��z�X����N$ݰ앫�;`pm`�| ���Da�rF1�"�-�U���Q݁��!8ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��~sj@��4B�-o��b����͟.O@��H'b6]��YjI]�8����c��H�q/�ɽ�*<e�7cϢA��z_'3�"�#F��8��5p���ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��S�"��[�#�Vxg�	h��(���!�(I�"j��5�{���	�����x�Y!"�#F��8S�B���@%����Z �jv�5�=���B���O�)��[��K�am@���h�n�gɽ�*<eɽ�*<eɽ�*<eɽ�*<e3la�nk�����N$��|�g�� k�kN�$�j������c�����|Gb��f	>���4�Qp?��y�ճ��:j���+���=a�^�ȕ����0��z#U�9�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e!��$и3�|��@S��ܦ���I��+r>[ؑ�#���vPt�8��5�쒈�R���%�^����<�e�/k�����tJe���״W�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w�7cϢA��[GK+��-��}%���Q�'Ws�t�����p�
�ӝE+<�u��y�ճ��:j���+���=a�^}4peOnɌ7X��q�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e!��$и3�p�������Ɛ�sg���ɒ(夜��=a�^:��鐗�ۄ��\��t\���OxO���<�e�/k����<�=�∿m���[̹ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w�7cϢA��[GK+����K�`�F����p������ O�bë�T�!���zN������%,!u�r�u^jP��:�(N�Ȟ��̸B��ຐ �R��;ɽ�*<eɽ�*<eɽ�*<e�VJUT��ȅV�)��w��Z�	/wx�ۻ�ٰ���˫��^���� Ĭ0w���W���̸B���Q�D@�ɽ�*<e�J�3fuza�^2�0�F�x�N8��ЎK�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����">̜��=a�^-��"�Kj���<���^R�:�`�<<�j!l���3)��q˃�6��Rbo� ���&ꬶ�R}�6'����_�,�\����]	M�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�E��!��~�]Sm�ʏY�u���)v%���©�U>�T@�͵�R}��_#��ц2�!��t��_�,�\��	(i{��y�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�E��!�R�M�"v�n�+�{_R��"�a��KlR41uz�s]eNN`ɽ�*<e��|P�f;��@�!���QFb�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��0'��n�v7����[��p����
��lz��4B�-旿�]��9�HF���,u�)�P��|P�f;��@�!݁��!8ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��0'��n@]�,��p���
��:�͟.O@��)v%���� O�bë�T�!���zN������P�O�_u^jP��:�[�-o�m�B����h�n�gɽ�*<eɽ�*<eɽ�*<e�VJUT���` �z�U; �C�a�jN<"�#F��8k�kN�$�Zŕ���EL*�����d<�xg��r��*�zN������P�O�_u^jP��:��D�!# ���"��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���` �z�U; �C�a�jN<�"vЅ\����ֿ74ı)v%����RC^��K�am@�&��r>�ɽ�*<e��|P� .=2��py<��֋���F��X
ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��0'��n���i�~R���*1��[��Ur�JFZŕ���E:(�\Ȝ��bb����Gk�w*o�Ё]-Ԗ����02v6cS&�*;��6�Geɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���` �z�U; �/�Ѭ��Na(�;�!�zS�e���QA��m��-��ڻ�y�ճ��vS+ё@�t�2M�����g�}��bWG��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e���>�(�J*/1Fu=S��;E�÷A����~��k�P˥V�7[c�a:~�9�[�P9��7�r�!��t��k�P˥-�{����:��Ҟ�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�E��!�{�����3�Q������}��a��v7�������z&AD*2�&I&ꬶ�R}�6'��ϗk�P˥���'B[t;�!�(I켚<dz�Uiɽ�*<eɽ�*<eɽ�*<e����n��r�E��!�{�����+)��S�*5V8��+ Z��F9R ��*/1Fu=S	/wx�ۻ����4�Qp?��y�ճ��vS+ё@�t�2M�����g�}}<��m�8��ЎK�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e���>�(�J�⧼��-�;YS�z(����<���^��?-h�j�v7����d+r9�N�����4�Qp?��y�ճ��vS+ё@�t�2M�c�A�`P���]	M�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e���>�(�J�⧼��-���D�do��ʏY�u���)v%�����>-����͵�R}��_#��ц2�!��t��R��+�����@�^�۳�EwW�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�E��!�t\����x����s�+X`NY̿��g.�I`�{d��T��zN������P�O�_��02v6c�p�s ���QFb�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���}�B-u��[��Ixۓ�S5�8x�XY��|P����MY��旿�]��9�HF���,u�)�P��|P�
a���aF.�;������m���[̹ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��0'��n���i�~R�lCi����K�`��F9R ��*/1Fu=So9�$�pD�H�q/�ɽ�*<e��|P�
a���aF.�[�-o�m�B����h�n�gɽ�*<eɽ�*<eɽ�*<e��0'��n���i�~R�lCi��"�#F��8k�kN�$�Zŕ���E[��Ixۓ������d<�xg��r��*�zN������P�O�_��02v6c�p�s ˃�6��Rb�<dz�Uiɽ�*<eɽ�*<eɽ�*<e�VJUT���` �z�U; љ.�;Xb>5xW�V8��+ Z��F9R ��*/1Fu=S���L��xg��r��*�zN������P�O�_��02v6c�ܠ
��d��!f�� �fɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���` �z�U; �:��*�$�EC���Z��e"��v7��������{%��ʶ��^��8�
���y��|P��Y�R�i�����BoܴW�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��0'��n���i�~R-���V-��}%���ƾYn��d�<g���p1	��S��`&ꬶ�R}�6'���ӿ�F��+ �Q� _9�传]�RH�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�)v%������
��Q�{���t�2M�'�'�N��q1�@"Z���y�ճ��0��hPz8�t�2M�� ���ƙ�8����c�>υU�%ߏɽ�*<eɽ�*<eɽ�*<eɽ�*<e���>�(�J�⧼��-�5�M���l���jX.Zŕ���E�,��\kb�ƚ�읻�y�ճ��vS+ё@�t�2M�� ���ƙ8�� �a����"��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e���>�(�J�⧼��-�W�7����JG5�td'���ֿ74ı)v%�����ھ�>j}�!�(I�o� ���&ꬶ�R}�6'���ӿ�F��+ ��>?��'��K�am@���h�n�gɽ�*<eɽ�*<eɽ�*<e����n��r�E��!�^4�LQ��"V��A|mk�kN�$�Zŕ���E�,��\kb�˃�6��Rbo� ���&ꬶ�R}�6'���41���) �)x5��;#tMɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�E��!�*v��U>t1jME���:��F9R ��*/1Fu=S�Gx5�th��b���cTk:�Р˵�t�2M�i?�����)	(i{��y�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e���>�(�J�⧼��-�'��~*�+�{_R��"�a���k��=�z�s]eNN`ɽ�*<e��|Pӛk�Oڴf�旿�]��Aв�2Gɽ�*<eɽ�*<eɽ�*<eɽ�*<e��0'��n�v7����샜/� �g��
��lz��02v6cBo
�=�L���ǅҸL�~bq�}pN<�W����02v6c�H1dȿ�݁��!8ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���` �z�U; y��8}v����
��:�͟.O@��)v%�������	�T�!���zN������P�O�_��02v6c�H1dȿ������d<�8��ЎK�ɽ�*<eɽ�*<eɽ�*<e�VJUT���` �z�U; y��8}v��}ɻ�&lc�̸B�����?-h�j�v7����=kpjg���m�B���&��r>�ɽ�*<e��|Pӛk�Oڴf���D�!# ���"��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��0'��n���i�~R+sF���5��"vЅ\����ֿ74ı)v%����f���GD�K�am@�&��r>�ɽ�*<e��|P�!M��chpy<��֋���F��X
ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��0'��n���i�~RH�7��[��Ur�JFZŕ���E5�%�A��bb����Gk�w*o�Ё]-Ԗ����02v6c�c�f�E����6�Geɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���` �z�U; �%�,K/�>�Na(�;�!�zS�e���QA��m��;t̴���y�ճ��vS+ё@�t�2M����^�'��bWG��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e���>�(�J*/1Fu=SU�ڻ9K�A����~�����>>�V�7[c�a:~�9�[�P9��7�r�!��t�����>>�-�{����:��Ҟ�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�E��!�=��� �3�Q������}��a��v7������,mɺ��AD*2�&I&ꬶ�R}�6'�������>>����'B[t;�!�(I켚<dz�Uiɽ�*<eɽ�*<eɽ�*<e����n��r�E��!�=��� �+)��S�*5V8��+ Z��F9R ��*/1Fu=S��(�4�1����4�Qp?��y�ճ��vS+ё@�t�2M����^�'}<��m�8��ЎK�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e���>�(�J�⧼��-��Ӻ0�������<���^��?-h�j�v7�����RE��и���4�Qp?��y�ճ��vS+ё@�t�2M�s��ĵ��&��]	M�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e���>�(�J�⧼��-���HB�x'�ʏY�u���)v%����2��c�x�͵�R}��_#��ц2�!��t�|�>��~����@�^�۳�EwW�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�E��!�	~q�j�mx����s�+X`NY̿�V�$�k��{d��T��zN������P�O�_��02v6c�1쀺T����QFb�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���}�B-u�Ö�YQy\�S5�8x�XY��|Pӡ�I;P��E旿�]��9�HF���,u�)�P��|Pӝqֺ|*��;������m���[̹ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��0'��n���i�~R�(�}��w��K�`��F9R ��*/1Fu=SKb���ÃH�q/�ɽ�*<e��|Pӝqֺ|*ӊ[�-o�m�B����h�n�gɽ�*<eɽ�*<eɽ�*<e��0'��n���i�~R�(�}��w"�#F��8k�kN�$�Zŕ���E��YQy\������d<�xg��r��*�zN������P�O�_��02v6c�1쀺T�˃�6��Rb�<dz�Uiɽ�*<eɽ�*<eɽ�*<e�VJUT���` �z�U; ��C�jli�>5xW�V8��+ Z��F9R ��*/1Fu=S{x�e�6�xg��r��*�zN������P�O�_��02v6c}i���Ҩ�!f�� �fɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���` �z�U; ��=�*��$�EC���Z��e"��v7����+��ެ.���ʶ��^��8�
���y��|P����������BoܴW�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��0'��n���i�~R< �Iـ�-��}%���ƾYn��d?���}1	��S��`&ꬶ�R}�6'��Ϸ Բ��+�Q� _9�传]�RH�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�)v%�����z4#R
�{���t�2M����_��pf1�@"Z���y�ճ��0��hPz8�t�2M����ܠ�Xџ8����c�>υU�%ߏɽ�*<eɽ�*<eɽ�*<eɽ�*<e���>�(�J�⧼��-�&�|�uu���jX.Zŕ���E�í�)��ƚ�읻�y�ճ��vS+ё@�t�2M����ܠ�X�8�� �a����"��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e���>�(�J�⧼��-����2ib�BG5�td'���ֿ74ı)v%���8p�!���!�(I�o� ���&ꬶ�R}�6'��Ϸ Բ��+��>?��'��K�am@���h�n�gɽ�*<eɽ�*<eɽ�*<e����n��r�E��!�i٥%��7"V��A|mk�kN�$�Zŕ���E�í�)��˃�6��Rbo� ���&ꬶ�R}�6'���s�(��|��) �)x5��;#tMɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�E��!��E�:�l��jME���:��F9R ��*/1Fu=SE�c�2-h��b���cTk:�Р˵�t�2M�Je�G%Ln	(i{��y�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e���>�(�J�⧼��-��lo!v%��+�{_R��"�a���ȟJ�gf�z�s]eNN`ɽ�*<e��|PӬyC�~|5旿�]��Aв�2Gɽ�*<eɽ�*<eɽ�*<eɽ�*<e��0'��n�v7����� J���m��
��lz��02v6c����P��L���ǅҸL�~bq�}pN<�W����02v6cP��
h݁��!8ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���` �z�U; )T��ׄHT���
��:�͟.O@��)v%�����!)=grT�!���zN������P�O�_��02v6cP��
h�����d<�8��ЎK�ɽ�*<eɽ�*<eɽ�*<e�VJUT���` �z�U; )T��ׄHT�}ɻ�&lc�̸B�����?-h�j�v7����A��*N2[�m�B���&��r>�ɽ�*<e��|PӬyC�~|5��D�!# ���"��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��0'��n���i�~R��ð����"vЅ\����ֿ74ı)v%���I�V������K�am@�&��r>�ɽ�*<e��|P�\ѯ
��?�py<��֋���F��X
ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��0'��n���i�~R�]mD��[��Ur�JFZŕ���Envh��J�bb����Gk�w*o�Ё]-Ԗ����02v6c#z�C-���6�Geɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���` �z�U; �/������Na(�;�!�zS�e���QA��mN�{��ٜ8��y�ճ��vS+ё@�t�2M�#����
1ͤ�bWG��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e���>�(�J*/1Fu=S�=�>H'A����~�L2�*<*S�V�7[c�a:~�9�[�P9��7�r�!��t�L2�*<*S�-�{����:��Ҟ�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�E��!�3�ge2�3�Q������}��a��v7����F �<�*AD*2�&I&ꬶ�R}�6'���L2�*<*S͋��'B[t;�!�(I켚<dz�Uiɽ�*<eɽ�*<eɽ�*<e����n��r�E��!�3�ge2�+)��S�*5V8��+ Z��F9R ��*/1Fu=S��D8QXz����4�Qp?��y�ճ��vS+ё@�t�2M�#����
1�}<��m�8��ЎK�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e���>�(�J�⧼��-�d�1��d���<���^��?-h�j�v7�������+��P���4�Qp?��y�ճ��vS+ё@�t�2M��� �O���]	M�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e���>�(�J`m�J�d ��p���آʏY�u���)v%���̻���
�5�쒈�R���%�^�n8��_`m�J�d3��� fT����8�:�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��|P�<W��4f%���Bo���F9R ��*/1Fu=Sm�O������y�ճ��vS+ё@�t�2M��� �Oत�bWG��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e���>�(�J*/1Fu=S�앫�;`p��F9R ��`m�J�dG:�}2 ˄ۄ��\��t\���OxOn8��_`m�J�d2�0g�2>��{���ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��|P�<W��4f%�;�������y��5}"�a��qQ	�K�BT�!���zN������P�O�_��02v6c�
�m���*�����d<�8��ЎK�ɽ�*<eɽ�*<eɽ�*<e�VJUT���` �z�U; NvX���_��}ɻ�&lc�̸B�����?-h�j�v7������htߧ�̸B���Q�D@�ɽ�*<e٫�,��9�5P,�>5xW�V8��+ Z�W�����ɽ�*<eɽ�*<eɽ�*<erL۪w�Ib�t�2M�]1�׮��}<��m�Ju9���ƾYn��d�C�&�J˃�6��Rbo� ���&ꬶ�R}�6'�����J������) �)x5��;#tMɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�E��!�
9.9T4�=jME���:��F9R ��*/1Fu=S�>fޅR�Mm`�| ��C4�X��E��!�Vnl�@�2��ʵ)n�{ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eeo9����02v6c�3�-݌O)ɠo>f�)v%����=(�%�ʥ1	��S��`&ꬶ�R}�6'�����J���׌Q� _9�传]�RH�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�)v%���+��ˏ�F�+ ���E��!�
9.9T4�=>�����m`�| ���Da�rF�E��!�Vnl�@�2�3�Q����M�tb�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eeo9����02v6c�3�-݌,�o��v+X`NY̿�r�e��aE����׃H�q/�ɽ�*<e��|P��lx���Ê[�-o�m�B����h�n�gɽ�*<eɽ�*<eɽ�*<e��0'��n���i�~R��B,Q���"�#F��8k�kN�$�Zŕ���ENRFb7H�"�#F��8S�B���@%����Zȩ�Ļ����i�~RڊQ��A8��"vЅ\�����}g�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e\T��}=l[��J������,�Ά�K�am@� 됰A�k��QA��mCZ�\:�(���4�Qp?��y�ճ��
�_�ڭWH��3�A�f<��T�;��.D#{?y���8�:�ɽ�*<eɽ�*<eɽ�*<e\�@?<���G:fGv��Y����#.cu,"y�zl>j�m�$Q��z�X e>oGn@al���ɡ���y�ճ���W7P�%����o=$W.����|c� k�k��L�����`�!f�� �fɽ�*<eɽ�*<eɽ�*<e�M,J����2���K,)e���.>��X�Bh�Wd��ٰ#s~^��n���l�ʶ�Pt�������q�ɚ G<��q��M�~���ySGQ��;ys2Ad ݰm�H/��+�ͼ�f���9TI��Vd?o9�ɽ�*<eɽ�*<eɽ�*<e[���g�Q����o=$W.����|������L�����`O)ɠo>fg�����6��o�����l!�ee1	��S��`&ꬶ�RQ�1	�|T�����)���W�X��<R|=-4Wj̼��Aв�2Gɽ�*<eɽ�*<e����n��rg�����6��o�������l�YZF�+ ����7�1��kC�������6�r&�����ڧ�P�7rV����ZMͿ���q�l�ʶ���u�[����h��_5��;#tMɽ�*<eɽ�*<eɽ�*<eɽ�*<e;���u�'�w�֬�ț����)�rj��+c5��)ϋ�2���K,)e���.>��X�Bh�W�	�y{I�7�͵�R}���JI#�a{�/%6�y
z'�w�֬��r}�<�P�p���[� ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rg�����6��o����h�rr�?A�O)ɠo>f��7�1��kC�������6�r�7Ց�X2͈��T�<����ZMͿ���q�l�ʶ���u�[��$�ss]d传]�RH�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��@�7�*T�����)�gUT�{<R|=-�z�`u�t�a�?�j��l�ʶ�Pt������$�ss]d:~�9�[�P�ǸX�e��/%6�y
z'�w�֬��r}�<�P�pzI�-�k��W�����ɽ�*<eɽ�*<eɽ�*<e����n��rg�����6��o����h�rr�?A����۾�t\dFK����f0%ڡ��u@G�ѥ䰾M^��i����m`�| �ɽ�*<e���{�}f$W.����|c� k�k��L�����`�!f�� �fɽ�*<eɽ�*<eɽ�*<e|�'B���ҫ�0�7�)e���.>��X�Bh�Wd��ٰ#s~^��n���l�ʶ���u�[���� �Y'��`v�ZP���܃$����~î�xa�-KB�i�Sd�~�fT�[V�`���S�)n%۳�EwW�ɽ�*<eɽ�*<eɽ�*<e�����ص�jU�.�S�9�tf���9TI�����7��G��S�'�w�֬����K��NF�ˀ����� �ɽ�*<e���'fLSx=��/��㟰��TM�B"�O�6a�s��ɽ�*<eɽ�*<eɽ�*<e���  I·]�찴�}0�@Z���ŗ߹������!����� �������jU�.�S�9�tf���9TI���.�NHm`�| �ɽ�*<eg�����6��o����a��רP��<1���F��X
ɽ�*<eɽ�*<eɽ�*<e�|�n����v2}&�PZ�n.{{�B�bty[[[��Ur�JF������Sx=��/��u@G�ѥ䰾M^� b��m`�| ����`�gg�����6��o����a��ר��))��W�����ɽ�*<eɽ�*<eɽ�*<e�|�n����v2}&�PZ�n.{{�B�bty[[-��}%��|�	R��-L�kC�������6�r�7Ց�X2͈��T�<����ZMͿ���q�l�ʶ���u�[����Ķ���U��bWG��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ص�jU�.�S�9�tf���9TI�I>/�4	���E�}X�v2}&�PZ�n.{{�B�bty[[�P�7rV����ZcP7�Ȯ��l�ʶ���u�[����Ķ���U�lƱOɽ�*<eɽ�*<eɽ�*<eɽ�*<e;���u�'�w�֬����K���GyE���EVWC�����{�}f$W.����|������%Y�g�E�wSj�F����ZЖ��ٿE
j���?�{�/z�p�^(]e��#J�����`��z#U�9�ɽ�*<eɽ�*<eɽ�*<e��@�7�*�-H嵰. �gUT�{<R|=-��X�Y6��H����&��v2}&�PZ�n.{{浐EÉ�1bb����G4�mJ�KZ�����)�ߙmit��Sd�~�fT�[V�`���S�)n%۳�EwW�ɽ�*<eɽ�*<e�VJUT���`Zʤ|�evA�^_p�x�S�9�tf���9TI�����7��G��S�'�w�֬���3��U��
NF�ˀ����� �ɽ�*<e��D�MA�^_p�x/��+�ͼ�f���9TI���.�NH�W�����ɽ�*<eɽ�*<e���  I·]�찴�}0�@Z���ŗ`�4�S��0!����� ��#�6KF5�-H嵰. �gUT�{<R|=-4Wj̼��9�HF���,ɽ�*<e�E�q�j��S�Y-�m`n��f��z�iU�}ɽ�*<eɽ�*<eɽ�*<ep<U˸����l�ʶ���u�[��M���p�iiͱH�R�#�6KF5�-H嵰. �gUT�{<R|=-}!�Lڜ<��q��M�~���ySG�,+�)c�B�2ƍ�zC�����y*8�����}۳�EwW�ɽ�*<eɽ�*<eɽ�*<e���  I·]�찴�}0�@Z���ŗ?��Sm
���~=���#�6KF5�-H嵰. �gUT�{<R|=-�n �u�HYz�s]eNN`ɽ�*<e�E�q�j��S�Y-�m`n�/"���S·�ۃRIɽ�*<eɽ�*<eɽ�*<e�:��MC��
j����M
��iͮp�^(]e����j�M�S5�8x�XY�E�q�j��S��8�ǧ/"���S�Ʒ2�v���䀒5k�,+�)c�B�2ƍ�zC�����y*��s$)?7`���kɽ�*<eɽ�*<eɽ�*<e���  I·]�찴�}0�@Z���ŗ?��Sm
�zI�-�k�5��)ϋ�}%^Y[�\V)e���.>��X�Bh�WJ8�-�3!L}�C2+�&ꬶ�RxP�Z�W揉ry�k����W�X��<R|=-��X�Y6����F��X
ɽ�*<eɽ�*<e����n��rn�>�B"�kC�������6�r&�����ڧ[��Ur�JF̵VA�T��B�2ƍ�zC�@Pek�#0�q�ɚ G<��q��M�~���ySGj�1���,S��c�P/��+�ͼ�f���9TI��Vd?o9�ɽ�*<eɽ�*<eɽ�*<e[���g�Q7��ɇ�F�$W.����|������L�����`O)ɠo>fg�����6��o����A'�
`���ϩ����Ȼ�y�ճ���W7P�%7��ɇ�F�$W.����|c� k�k��L�����`���QFb�ɽ�*<eɽ�*<eɽ�*<eVӥRysL_��v������D�Oȝ��Iy��0F�+ ��n�>�B"�kC�������6�r&�����ڧ�P�7rV����ZMͿ���q�l�ʶ���u�[��G1~l��҆��]	M�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e;���u�'�w�֬���AV�n��j�"X�ʏY�u��n�>�B"�kC�������6�r�7Ց�X2l���ɡ���y�ճ���FʄL�)�]�찴�}0�@Z���ŗ AM��jt���[� ɽ�*<eɽ�*<eɽ�*<eɽ�*<eVӥRysL_��v������D�OȝڙcS����O)ɠo>fn�>�B"�kC�������6�r�7Ց�X2͈��T�<����ZMͿ���q�l�ʶ���u�[��G1~l��҆��bWG��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�iƅ��ry�k��gUT�{<R|=-�z�`u�t�a�?�j��l�ʶ���u�[��B�����1�@"Z���y�ճ��u�@T�t��]�찴�}0�@Z���ŗ AM��jtzI�-�k��W�����ɽ�*<eɽ�*<eɽ�*<eVӥRysL_��v������D�OȝڙcS�������۾�t\��Z0B��)�xoĪ��u@G�ѥ䰾M^��i����m`�| �ɽ�*<e|2w�e�Q��kC����^��N2�{�&�����ڧ7R��ɽ�*<eɽ�*<eɽ�*<e|�'B����I�\�m�ʽ�ʾ�ց[V�`��zǙ�7��&u
1�F�]�찴�}0�@Z���ŗ�?Zd��&��ؒ��y�ճ���QGK�z	RIꐦO�j$W.����|c� k�k��L�����`��6�Geɽ�*<eɽ�*<eɽ�*<e�M,J���܁����=�)e���.>��X�Bh�W�0���Ѓ�j�ğ %D�v2}&�PZ�n.{{M���=s�i��g��Z�����Ť2��9�|�����=����3e�X�Bh�W.����T�3·�ۃRIɽ�*<eɽ�*<e,4���?w�E�q�j��S�{�/������N�U��!�L?7Ƌ�I�\�m�ʽ�ʾ�ց[V�`��,\�8� 'z:~�9�[�P&ꬶ�R\���d!2'�w�֬�ȇ��nD�NJ��� ��z#U�9�ɽ�*<eɽ�*<eɽ�*<e����n��rg�����6��o����}K��'�P��<1��!�"
��u�I�\�m�ʽ�ʾ�ց[V�`���>Q�����5�쒈�Kv@�tsQ���g����v������D�Oȝ��QL�~P��6�Geɽ�*<eɽ�*<eɽ�*<e,4���?w�E�q�j��S�ͼW�S0cnW8���2D�5�O��I�\�m�ʽ�ʾ�ց[V�`���>��h�
1	��S��`&ꬶ�R\���d!2'�w�֬�ȇ��nD�<�䴗�.��7X��q�ɽ�*<eɽ�*<eɽ�*<e����n��r|2w�e�Q��kC�������6�r�7Ց�X2�ѥ������G��S�'�w�֬�ȇ��nD�x*0��ۄ��\��t3>1]Q-y���g����v������D�Oȝ��QL�~P;*[��Fɽ�*<eɽ�*<eɽ�*<e,4���?w�E�q�j��S�ͼW�S0c�N�y��^Cb��D8>�u��	�d��M
��iͮp�^(]e����j�M�%E5fT��zN�����1稆���%��+ v���Sd�~�fT�[V�`��zǙ�7�5��;#tMɽ�*<eɽ�*<e�VJUT������9f?��;�T�S�9�tf���9TI��~-y7�f-�ž嫆v������D�Oȝ����u�^�5�쒈�Kv@�tsQW|9��\�ڇ��C������3e�X�Bh�W�0���Ѓ�x`һaB�ɽ�*<eɽ�*<e,4���?w��Z0B��n�Rd%���u@G�TM�B"�O&0�w��̵VA�T��B�2ƍ�zC�y;�R���_<��D��z�s]eNN`ɽ�*<e��Z0B��n�Rd%���㟰��TM�B"�O�6a�s��ɽ�*<eɽ�*<eɽ�*<ep<U˸����l�ʶ���u�[������F��.���Ȁ���,d�?���;�T�S�9�tf���9TI���.�NHm`�| �ɽ�*<eg�����6��o�����B-�>�P��<1���F��X
ɽ�*<eɽ�*<eɽ�*<e�|�n����v2}&�PZ�n.{{'��{�k[��Ur�JF��,d�?���;�T�S�9�tf���9TI'�09k� ���ʶ��^ͮ��f�?�E�q�j��S�5��ȺTanW8���x`һaB�ɽ�*<eɽ�*<eɽ�*<ep<U˸����l�ʶ���u�[��R�\����� 
�KO���,d�?���;�T�S�9�tf���9TI�;�Y��##m`�| �ɽ�*<eg�����6��o�����B-�>��d��2��.Aв�2Gɽ�*<eɽ�*<eɽ�*<e|�'B�����+ v����ʾ�ց[V�`��G	�ģ�BF�+ ��g�����6��o����>��B��;��d��2��.9�HF���,�-� ����E�q�j��S�5��ȺTa�N�y��^C��N�mp�ɽ�*<eɽ�*<eɽ�*<ep<U˸����l�ʶ���u�[��R�\������g}��nAX�
�j�3Ɖ�D��0L�gUT�{<R|=-�;�����}��
΄ɽ�*<e�@������Ժ��h�/��+�ͼ�f���9TI��~-y7�W�����ɽ�*<eɽ�*<e[���g�Q�ϝO�}�$W.����|������L�����`0�ۧ��5��E�q�j��S�
�Y�w�)]gpSPJeX��ʶ��^ͮ��f�?��Z0B��N'�������㟰��TM�B"�O��5_m��ɽ�*<eɽ�*<eɽ�*<e�:��MC��|m9T�g�R�M
��iͮp�^(]e��A ��%@�����c]�찴�}0�@Z���ŗ��e�h�I͟ܜ��������ZЖ��ٿE|m9T�g�R?�{�/z�p�^(]e��C�]�Nf�݌7X��q�ɽ�*<eɽ�*<eɽ�*<e;���u�'�w�֬��-��?H!3@��=)����
�,��,�ϝO�}�$W.����|������L�����`L���ǅҀzN������7l&��F��v2}&�PZ�n.{{~25!��`7R��ɽ�*<eɽ�*<eɽ�*<e�VJUT��� �H4%B�2ƍ�zC1aXW�b�ف�h��_����G8�ϝO�}�$W.����|������%Y�g�E��`v�ZP���܃$���80��k ���l�ʶ���u�[��|_�Nſ	(i{��y�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e;���u�'�w�֬��-��?H!3(��{�Ը�x-L
��ϝO�}�$W.����|������%Y�g�E��{d��T��zN������7l&��F��v2}&�PZ�n.{{~25!��`b:n\��ɽ�*<eɽ�*<eɽ�*<e�VJUT������9f?��Ժ��h��S�9�tf���9TI�I>/�4	���E�}X�v2}&�PZ�n.{{pH�#ʷ�P�7rV����ZcP7�Ȯ��l�ʶ���u�[��|_�Nſ�lƱOɽ�*<eɽ�*<eɽ�*<eɽ�*<e;���u�'�w�֬��-��?H!3�GyE���EVWC����3����kC�������6�r�7Ց�X2�[�S�BtM��y�ճ���W7P�%(�2Y�ǫ$W.����|c� k�k��L�����`�!f�� �fɽ�*<eɽ�*<eɽ�*<e�M,J���ܕpᓖC�)e���.>��X�Bh�Wd��ٰ#s~^��n���l�ʶ���u�[���ƴh	L�`v�ZP���܃$����~î�xa�;i���`C>?�{�/z�p�^(]e��A ��%����8�:�ɽ�*<eɽ�*<eɽ�*<e�iƅ�����N�B�gUT�{<R|=-}��&�rS�f-�ž嫆v������D�Oȝ�%6��1	��S��`&ꬶ�RxP�Z�W揗���N�B���W�X��<R|=-4Wj̼��Aв�2Gɽ�*<eɽ�*<e����n��rg�����6��o�����
m���U��&�}5��)ϋ��pᓖC�)e���.>��X�Bh�W.����T�3�Ʒ2�v�ɽ�*<e@82�����B�2ƍ�zC�c���b��h��_5��;#tMɽ�*<eɽ�*<eɽ�*<e���  I·]�찴�}0�@Z���ŗ//l���w)�rj��+c5��)ϋ��pᓖC�)e���.>��X�Bh�W�	�y{I�7�͵�R}���JI#�a{�/%6�y
z'�w�֬��n�r#�O1j�����0����8�:�ɽ�*<eɽ�*<eɽ�*<e����n��rg�����6��o�����I&�s���))�5��)ϋ��pᓖC�)e���.>��X�Bh�WC'�K��w���� �ɽ�*<e@82�����B�2ƍ�zC�c���b$�ss]d传]�RH�ɽ�*<eɽ�*<eɽ�*<e[���g�Q(�2Y�ǫ$W.����|������%Y�g�E��.���Ȁ�̵VA�T��B�2ƍ�zCw	z9���$�ss]d:~�9�[�P�ǸX�e��/%6�y
z'�w�֬��n�r#�O1{M)����h3a�̌Kɽ�*<eɽ�*<eɽ�*<e����n��rg�����6��o�����I&�s�O4����UZ�Ԯa���u�6�f�3��ʾ�ց[V�`�����@��=����Z�����Ť2��9�|H���5������3e�X�Bh�Wd��ٰ#s�z�iU�}ɽ�*<eɽ�*<e,4���?w��Z0B��2h�L�&�_��u@G�TM�B"�Ol>j�m���G��S�'�w�֬��2:���f~�)��C��͵�R}���JI#�a{aV�CF�[�
��S�V���W�X��<R|=-}��&�rS�W�����ɽ�*<eɽ�*<e����n��r�/�ӄi�4�kC�������6�r&�����ڧ-��}%���E�q�j��S��^�ϤW���KS�m`�| �ɽ�*<e�/�ӄi�4�kC����^��N2�{�&�����ڧb:n\��ɽ�*<eɽ�*<eɽ�*<e�|�n����v2}&�PZ�n.{{"�EB6gW6S5�8x�XY��Z0B��2h�L�&�_��u@G�TM�B"�OM'6/�`��y�ճ��kwO�&뿃]�찴�}0�@Z���ŗ��qy�6�)�rj��+c�W�����ɽ�*<eɽ�*<eɽ�*<eVӥRysL_��v������D�Oȝ0+H,�"k�0�ۧ��5���Z0B��2h�L�&�_��u@G�ѥ䰾M^� b��m`�| ����`�gg�����6��o����-V�P�����))��W�����ɽ�*<eɽ�*<eɽ�*<e�|�n����v2}&�PZ�n.{{;��v�_-��}%����Z0B��2h�L�&�_��u@G�ѥ䰾M^r/�0!�$���y�ճ��kwO�&뿃]�찴�}0�@Z���ŗ��qy�6�U��&�}�W�����ɽ�*<eɽ�*<eɽ�*<e�M,J����H���5�)e���.>��X�Bh�W��.����A��m.x�^]�찴�}0�@Z���ŗU5���
�U��&�}m`�| ���"�v�h�g�����6��o����-V�P���O4����U�Q���)8�ɽ�*<eɽ�*<eɽ�*<e�|�n����v2}&�PZ�n.{{;��v�_݀���b���,d�?���f���S�9�tf���9TI�&!�r8�s��}v�h�ɽ�*<e��Z0B�����V�����㟰��TM�B"�OX P��>d}ɽ�*<eɽ�*<eɽ�*<e�:��MC�٩`���$���M
��iͮp�^(]e��#J�����`�ʏY�u��g�����6��o�����'�Ad�Ȧ)�rj��+cm`�| ����`�g��?��B��kC����^��N2�{�&�����ڧ�S�P'qɽ�*<eɽ�*<eɽ�*<e|�'B���;	��7�8��ʾ�ց[V�`���S�)n%��oB���l�ʶ���u�[�������S�{d��T��zN�����1稆���%;	��7�8�Sd�~�fT�[V�`��,\�8� 'z传]�RH�ɽ�*<eɽ�*<e�VJUT��� �H4%B�2ƍ�zC�;t�Ս��^Ii6Q�,��/�`���$���M
��iͮp�^(]e��C�]�Nf��ۄ��\��tZ�����ŕ~�}������v������D�Oȝ�)��>�!f�� �fɽ�*<eɽ�*<eɽ�*<e,4���?w�E�q�j��S��8
���-��f�8�̣*��ة`���$���M
��iͮp�^(]e����j�M�bb����G4�mJ�K�YU�@N���v2}&�PZ�n.{{��;����S�P'qɽ�*<eɽ�*<eɽ�*<e�VJUT��� �H4%B�2ƍ�zC�;t�Ս8�����}=�n\��{J�`���$���M
��iͮp�^(]e����j�M��i��g��Z�����ŕ~�}������v������D�Oȝ�)��>���QFb�ɽ�*<eɽ�*<eɽ�*<e,4���?w��Z0B�����V�����u@G�ѥ䰾M^�������f-�ž嫆v������D�Oȝ�����, ?L���ǅҰ#�L��פ���Ԡ�T�v2}&�PZ�n.{{��;�����g���;�ɽ�*<eɽ�*<eɽ�*<e�VJUT��� �H4%B�2ƍ�zC�;t�Ս��s$)`PF�ꇜ��s7�}��$W.����|������%Y�g�E�wSj�F����ZЖ��ٿEm��3+� �?�{�/z�p�^(]e��#J�����`��z#U�9�ɽ�*<eɽ�*<eɽ�*<e�iƅ�C�6�vm��gUT�{<R|=-��X�Y6��H����&��v2}&�PZ�n.{{�q�"��\fbb����G4�mJ�KZ�����@w������Sd�~�fT�[V�`���S�)n%۳�EwW�ɽ�*<eɽ�*<e�VJUT������9f?(�&���S�9�tf���9TI�����7��G��S�'�w�֬���D;�k�NF�ˀ����� �ɽ�*<e�@����(�&��/��+�ͼ�f���9TI���.�NH�W�����ɽ�*<eɽ�*<e���  I·]�찴�}0�@Z���ŗ+�_X��!�!����� �X�
�j�3C�6�vm��gUT�{<R|=-4Wj̼��9�HF���,ɽ�*<e�E�q�j��S����k3��f��z�iU�}ɽ�*<eɽ�*<eɽ�*<ep<U˸����l�ʶ���u�[��I�pù��iiͱH�RX�
�j�3C�6�vm��gUT�{<R|=-}!�Lڜ<��q��M�~���ySG�,+�)c�B�2ƍ�zC>��@��8�8�����}۳�EwW�ɽ�*<eɽ�*<eɽ�*<e���  I·]�찴�}0�@Z���ŗ���:�-��~=���X�
�j�3C�6�vm��gUT�{<R|=-�n �u�HYz�s]eNN`ɽ�*<e�E�q�j��S����k3�/"���S·�ۃRIɽ�*<eɽ�*<eɽ�*<e�:��MC��m��3+� ��M
��iͮp�^(]e����j�M�S5�8x�XY�E�q�j��S���>�|��M�/"���S�Ʒ2�v���䀒5k�,+�)c�B�2ƍ�zC>��@��8���s$)?7`���kɽ�*<eɽ�*<eɽ�*<e���  I·]�찴�}0�@Z���ŗ���:�-zI�-�k�5��)ϋ� �D�O�h>)e���.>��X�Bh�WJ8�-�3!L}�C2+�&ꬶ�RqZKǅ�u'a���g�_��㟰��TM�B"�OX P��>d}ɽ�*<eɽ�*<eɽ�*<e����n��r�c�i�#J�M
��iͮp�^(]e��#J�����`�ʏY�u��g�����6��o�����.ץ/:��)�rj��+cm`�| ����`�g�c�i�#J?�{�/z�p�^(]e��A ��%����8�:�ɽ�*<eɽ�*<eɽ�*<e|�'B���׷�����0�gUT�{<R|=-}��&�rS�f-�ž嫆v���@�/���H ���P�1	��S��`&ꬶ�RqZKǅ�u'a���g�_��㟰��TM�B"�O�6a�s��ɽ�*<eɽ�*<eɽ�*<e����n��rg�����6��o�����.ץ/:��U��&�}5��)ϋ���;��Y��S�9�tf���9TI���.�NHm`�| �ɽ�*<eg�����6��o����1�ƚ��P��<1���F��X
ɽ�*<eɽ�*<eɽ�*<e�|�n����v2}&�PZ�n.{{��Z[)�[��Ur�JF�w��nR>��kC�������6�r�7Ց�X2l���ɡ���y�ճ���FʄL�)�]�찴�}0�@Z���ŗ��ݐ�1���[� ɽ�*<eɽ�*<eɽ�*<eɽ�*<eVӥRysL_��v���@�/����#��Iװ�O)ɠo>f�c�i�#J�M
��iͮp�^(]e����j�M��i��g��Z�����ŕ~�}������v���@�/�������ys/���QFb�ɽ�*<eɽ�*<eɽ�*<e,4���?w�+T��u0�$W.����|������%Y�g�E��.���Ȁ�̵VA�T��B�2ƍ�zCX��0/��$�ss]d:~�9�[�P�ǸX�e��/%6�y
z'�w�֬�Ț�/�� ��{M)����h3a�̌Kɽ�*<eɽ�*<eɽ�*<e����n��rg�����6��o������A-Tq�O4����UZ�Ԯa��׷�����0�gUT�{<R|=-�;�����@�{��Uⳮ3f�d
��v�g˨�&�;���`j�{=�}\��8B`}�FW,P���� ��蠀�&�Ī;��ɽ�*<eL�@t�Z�sȩ�h�<L8���5V��ɽ�*<eɽ�*<e-&�
:lݲ|PZ��9ԁQ�onv>�v2DaZqOɽ�*<e}���5�lt���/B���5���ɽ�*<eWO`&뼪f��+O��yu")�
B����]iLɽ�*<e�A����׏��w��C����L�N�����]iLN9�-(�/��!���7�%ܒ��5H�ɽ�*<eɽ�*<e�%�G��,���,	F��ݏ�ɽ�*<e�tO�4�!���7�%F�$��]!�#lѥ��X��Ɍw\�d��JęS�?�4�AT͗|Gn��(i��;k.n��U�ۄ���!���7�%��<2a'K̐I�rɽ�*<ed��Ję ���ga+D��'���ɽ�*<e��U�ۄ���!���7�%����jCORuI��<ɽ�*<e�%�G��"�! �^О�UC
��ɽ�*<e�tO�4�!���7�%fKˍʔ��	kU�f�Zɽ�*<ed��Ję�,���,���=��Z���s��[��U�ۄ����S��$�w�&��y�2 �9bA��ɽ�*<e�dtD<]�<�AP����k ��y$���>�|��
�tO�4��S��$�ws�m]��ȋ,�F��f�g6�S('�d��Ję�#�כnp���4�MS5�w:ɂ���s�EŖڿ=���ھ��:^��ġ��N���d��Ję©�yJ��j�=�+1�Vn���3��U�ۄ����S��$�wK��G�>@V�d!��X{t85�T-�$��8����\���ֻ'r�f�'��Sb�&9��̹尮l;�DhY��F�ɽ�*<e1? ��6�+t�c�K�]��s�kɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<eɽ�*<e-��fΡ��k��4t�pԖ�����Mhɽ�*<e�Y��2�K+��Qݓ˟s4�)�_π ����������'�e����ǄQ�]�Q�Mɽ�*<eɽ�*<e�����ɽ�*<evS+ё@�˴qZ5�g�}4"{t��HN�E���>Է4�Y�3�9��F�t�e�Q��8��y	&-l���P|P�퍓�rlV)iz������$���
���2�h
�K=4VӥRysL_ �1J�`���'t,�|n@��.�oԣ�;�d ��Ol��
��w_�}�X"nɽ�*<e�������Br(�&G!1���s�D�<@m̞���&m(��ϑi���8x���`�U�Q	76
m�"�x�\�uɽ�*<eɽ�*<eɽ�*<e��"�m҂B�1ci��)�<�;ɽ�*<e@�j/�j��ڭWH��EZ)eb?S�)��ש0��y�;Xz�����phl���q|���AQ�OsJɽ�*<eNM{9q��ɽ�*<eɽ�*<e�H��g�h�Q���:q����d�ɽ�*<e@�j/�j��ڭWH��EZ)eb?S�)��ש0��y�;Xz�����phl���q|���˟M�o}Q�]�Q�MNM{9q��ɽ�*<eɽ�*<e��vVK�`���;�	E\��М}��(H��u�6��/���%�\���ֻ'r�f�'��Sb�&9�����ڎXJ��&�+{����W&[��O�>�5��2��AqzY[v�_�ɽ�*<eɽ�*<e+�n�/�G��rq��&��sQ��~=��O��b2�M/��J@�j/�j��ڭWH��EZ)eb?S�)��ש0��y�;Xz�����phl���q|����f>;�݃����h��,K�%-
+[ɽ�*<eɽ�*<e�H��g澁_d�Ǹ��#��6*+�'�(.%�,aކ���jq�/���%�\���ֻ'r�f�'��Sb�&9�����ڎXJ��&�+{����W&[�a� ��^�$�c>y�DY[v�_�ɽ�*<eɽ�*<e+�n�/�G���g�#w�O!#Y��y�P����g��������Y�3�9��F�t�e�Q��8��y	&-l���P|P�퍓�rlV)iz������$��P�6;7}�&ZReX�ҝ[��R�ɽ�*<eɽ�*<e!�T9�u�P�+H�"hb��e�dB�$Dɽ�*<e��@�� ���q|���mVW��c�=��[�sr�G�^6,v��n��g���݇\��D��M�N�����n��rɽ�*<eɽ�*<eɽ�*<e��DO�y4�a����"G��0�@��ɽ�*<e@�j/�j��ڭWH��EZ)eb?S�)��ש0��y�;Xz�����phl���q|���U���g(ɽ�*<eNM{9q��ɽ�*<eɽ�*<e?������|�ޒ�j\S���Γ1��#�s@�j/�j��ڭWH��EZ)eb?S�)��ש0��y�;Xz�����phl���q|����>��܎�E#L�@���NM{9q��ɽ�*<eɽ�*<e��Ԫ�N��Lj}��i�S]�O{ݱ��
���2ɽ�*<e�Y�3�9��F�t�e�c���L)�/'~_�~Nɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R��E�q�j�����0n@��.�oԣ�;�d ���Y�n���(H��u�6�ɽ�*<e�������i�OϿY�M�L>�;>cc��R��Mbɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<eɽ�*<eɽ�*<e0��葠�Q���Д4��V�3yn�3y֜�V����/���%�\���ֻ'�ȡ�X0���b\	y`��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<eɽ�*<e+�n�/�G���g�#w!��zi"���IPd��Qɽ�*<e�Y�3�9��F�t�e�'l�����d�h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<eɽ�*<e!�T9�G�S$
�п�P�6;7}49�iv (�Y�3�9��F�t�e�'l�����dw�	�6�cɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<eɽ�*<e!�T9�u�P�+H�"Sv(a�iP��%e�܉�j�<�U�q��@�� ���q|���/���?���AE
!�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<eɽ�*<eɽ�*<e7[��İ��f�Ӗ�F>�8��O6�QWk�HZ�ɽ�*<eS*��j��ΗCf�|�"���y��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<eɽ�*<eɽ�*<e�]Ӟv��H�p^|��]`�ɽ�*<e�����+���G:fGv��LQ{D��y�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<��ɽ�*<eɽ�*<e��r���
�JP$�I��u+��(W����sp�ɽ�*<e��Ԗ�ejɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e��p�^���Lc ��9t����� 3��;x�J�u�CK�U�}�q26�\�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e��=�wYh�ǵ��Љ�>>z�c��<��iP��[P-&J�� ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e��p�^���Lc ��9t����_�av"	;��%������z:�-q26�\�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e��=�wYh�ǵ�t:�󫓔ɽ�*<eɽ�*<e-&J�� ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e��p�^���Lc ��9t���ɕ?kV7�(T�F(�œ��z:�-q26�\�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e��=�wYh�ǵ���c{Qb�!�Z��ɽ�*<e�����l�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e��p�^���Lc ��9t�����T-��|�ɽ�*<e���z:�-��t$��oɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e��=�wYh�ǵ����#�H˥�j����N0ɽ�*<e�����E-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e��p�^���Lc ��9t���\#����r�ɽ�*<e������ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e��=�wYh�ǵ공�h�Ɔ�L{���V݅Ϗm�/
-&J�� ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e��p�^���Lc ��9t������(�-����)P�hx�-��m�[$ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e��=�wY�@o��W������&�5G���0��Jf�x�\("mVW��c�=H\�p�θ��Ɯ�h�[�Z�~�qe'%��@�|)��t���ɽ�*<e�/���%�ȩ�h�<L8���5V��ɽ�*<eɽ�*<eL�@t�Z�sv/G�ˀ��uۨ�T���]iLɽ�*<eL�@t�Z�sȩ�h�<L8��=HI~��a�l��ɽ�*<e�+ �0��0�{��NȈUP�h~��LZ\8��.��ɽ�*<e�tO�4s�EŖڿUP�h~��LZ\8��.��ɽ�*<eWO`&뼪f��+O��yu")�
B����]iLɽ�*<e-&�
:lݲf��+O��s�m]��ȋ��ϋ8z��ɽ�*<e�I*{_���"�}�H��ڳ�/��I�U�Z�ɽ�*<e�.���)V�T(�<7�l��FO�T��
��i�ɽ�*<ed��Ję"�! �^О�UC
��ɽ�*<eɽ�*<e�ߐuX�q��]6�*�z�&�=�34ɽ�*<e�/���%󬧁��ȉ�iOD�ɕ�U�_rw���+ɽ�*<e-��)ӕyL��P�a��$���$t�_rw���+ɽ�*<e��U�ۄ����S��$�w�&��y�2 �9bA��ɽ�*<eWO`&뼪嬷b
�{F���Y�ĀS��ɟ��ɽ�*<e7�3]N|�d���7{�n�5Ǔ��G|3k.sb}ɽ�*<e�.���)V��������8<NDD�{O��8{�U7-{�$0�d��Ję��I}�8<NDD�{O��8{�U7-{�$0��ߐuX�q�t7I�鄂|#e�;��JH5c�҃�pBT�7��t擱���I_��Ú�ȩ�F�(Uo��f�,+��a�����}0�{��NȈ���R���]В����E���bT�>�tO�4��S��$�w�	��?�K(В����E���bT�>�U��h����R��z�{dG`��Z"c���Y��ɽ�*<e7�3]N|���� &��U��GBM�J=P�P9Qɽ�*<erP/�ۻ�dFK��/��J��o�u�����` 0��%rɽ�*<eɽ�*<eǋ'H)�@w����a���h
�K=4ɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<eɽ�*<e-��fΡ��k��4t�pԖ�����Mhɽ�*<e�Y��2�K+��Qݓ˟s4�)�_π ����������'�e����Ǆ,K�%-
+[ɽ�*<eɽ�*<e����F���� �\����8��#�˴��56$����sb����o=$W.����|txG�z��h'~_�~Nɽ�*<e���  I·P|P�퍓�rlV)i��F}�~RΔm��ڡ^J�h��J�EL�cm�wo�	h�[�,��T"��T�����)�堒�c��[�eonDS2��Y5��ɽ�*<e�����ɽ�*<eɽ�*<e�LOG۳=���f���B}�k���"�l��Z=�ɽ�*<emD�ْ�Ad ݰm�H2� ���TD�>蔽iɽ�*<e�VJUT���?�(<��ɽ�*<eɽ�*<e�bv�t>W�|m:�w�Ef�af�w�ɽ�*<e�,��T"��T�����)�堒�c�k;c���xɽ�*<eɽ�*<e�����ɽ�*<eɽ�*<e��r�Ϻ�0�7��R���7��$`љR��Y��2�K+A�O�����`�f ��{I����!����$e6ɽ�*<eNM{9q��ɽ�*<eɽ�*<eZi��LύE��9�����fQ�΀��P�6;7}�~�p[�3�Y��2�K+A�O�����`�f ��{�f>;�݃����h��Q�]�Q�MNM{9q��ɽ�*<eɽ�*<e!�T9���z�IYLyǺ �v�$V�3yn�3y֜�V���$����sb����o=$W.����|Fɱ�˕���2���}�ɽ�*<ex�\�uɽ�*<eɽ�*<e+�n�/�G���g�#w�O!#Y��y�P����g�������X��~?�W#��}��N?�{�/z�eg�/��y�����ɽ�*<eY[v�_�ɽ�*<eɽ�*<e�H��g澚c����|m:�w�E^|��]`�ɽ�*<e�,��T"��T�����)�堒�c�i���!�)��&ZReX�ɽ�*<e�����ɽ�*<eɽ�*<e��r���
�JP$��)3LQuq�DhY��F�ɽ�*<eO��'��f0%ڡ��8�z4ؓ���+4�ɽ�*<e,4���?wɽ�*<eɽ�*<eɽ�*<e	���j��7��9�G,�IM�+�I���>Է4mD�ْ�Ad ݰm�H94���i�Lj}��	�q��IX;�VJUT���?�(<��ɽ�*<eɽ�*<e���|���(zSȢ�|�RhꭣLš�	"�$ɽ�*<emD�ْ�������d��}�o���ɽ�*<eɽ�*<e�VJUT���\�ȱ���P��o��@G,6�`|yiglW�yi�S]�O{ݿ�P�6;7}49�iv (X��~?�W#��}��N�hM'��IN�\U�>:�ɽ�*<eɽ�*<eY[v�_�ɽ�*<eɽ�*<e�H��g澚c�����8��O6�QWk�HZ�ɽ�*<e�^1�?q�-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\U9��8P���)�<�;ɽ�*<e�/���%��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc ��9t���i���!�)�49�iv (������ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%�)0�/ئ�C�Ȩ_�����2�H���A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%���������DC�M�f��E�-MZ�F�Aܘ���E���m'Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���mg��gT�wJ�EL�cm�wo�	h�[i=�Z ���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��=�wYh�ǵ�7����h=aކ���jqɽ�*<e�����l�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡN��Y�T�P�6;7}�~�p[�3�	���t�nj�'%萚 tɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�fmC���|��9���wo�	h�[S�;��$�Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\U9��8P�q����dל��g�#w�lm�l1�b�h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc ��9t�����p��,ɽ�*<e������ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%� �G�\�<��;�sɽ�*<e��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%���������DC�Mx�-8��kɽ�*<ea�磅"��Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���m��G�I�9��T-��|�ɽ�*<e��{��Q�h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��=�wYh�ǵ�敥�2��t:���y��Vɽ�*<e�����l�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡN��Y�T�ͤ����ly֜�V�������pɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�f'����c���ڇ
�܎[ɽ�*<e�^1�?q�-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\U9��8P�5�ר��M^��i�?�/���%���U�?��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc �P�~Y���p)2���@�h2uv�%��k�{4ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%$-͇����L{���V݅Ϗm�/
UXec��
ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%������R
�CI���$�$�w�'�����j){rM
���אSb�&9��b��i���sX!�*����)A ˯nkB�J�tx�E�Bxɽ�*<e=���DХ��S��$�wP�.a7)�ɽ�*<eɽ�*<e[a�?~��s�EŖڿ�K[�k�ɽ�*<eɽ�*<e[a�?~����S��$�ws�m]��ȋ��ϋ8z��ɽ�*<eݵYi�|PZ��9ԁl]:G�&C�L5��eɽ�*<e�
���Wϓ��D��C��l]:G�&C�L5��eɽ�*<e�!�o�5���e�q>$��ޘ ~��fɽ�*<eɽ�*<e^iB�j��� UI�!n�5Ǔ��G�tx�E�Bxɽ�*<e$Q0��0���� <�n�S����{ɽ�*<eɽ�*<e�ߐuX�q�&2}��$R�����aO�!��/���%󬧁��ȉ�iXv���VF�@��C ��ɽ�*<e-��)ӕyL��P�a��B/Pb��|�\��7��ɽ�*<e��U�ۄ���!���7�%fKˍʔ��	kU�f�Zɽ�*<e�U��h���Lw��c����^pl	kU�f�Zɽ�*<e7�3]N|�R�RN@����R5�+ұ�i�A[�%ѯɽ�*<e�!�o�5���� ��蠀����N�!?�iRiɽ�*<ed��Ję��NYu._Zf3�����S��ɟ��ɽ�*<e�ߐuX�q�l���]6��쵪9s�����	֭U����[�����ȉ�il���]6��쵪9s�����	��z��X��0�{��NȈf����u�J�[�[�d���7�y��|�{�V`Z]�������>X����ݞ��d/�)�+j�9)@À)U�~\�80R���<y?�Bd:�6�}Zɽ�*<e�
���Wϓ$0D�7����uĥN�Bd:�6�}Zɽ�*<e�.���)VG%�"�}Ɗ��G�o��J=P�P9Qɽ�*<ed��Ję�	�ګ���+��n�X�J%�Y��ɽ�*<es�HB	�k�F{N.JIK�vv��O�ơ���a'ѳ��w��ɽ�*<eɽ�*<e��=!��(2��p�ɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<��ɽ�*<e:j���+�oaf�	��,��/�=X]ɽ�*<eɽ�*<emD�ْ�dh89QN��hz�;3��PY���F��
�W���[�&���2�%?�(<��ɽ�*<e��_��l���<I}���G�I�9w��\��ɽ�*<e[��ղ�f�!��QE���堒�c�)u/��L�<Q�]�Q�Mɽ�*<eVӥRysL_ �1J�`���u@�:4j�ק�	��� 4���:o�W��JW����sp��/���%󬷌�{�}f$W.����|Y�<d�2!#	76
m�"�ɽ�*<e����n��rɽ�*<eɽ�*<eɽ�*<e��"�m҂B�1ci��)�<�;ɽ�*<e$����sb�F{N.J?�{�/z�&�d}�=cUQ�]�Q�Mɽ�*<ex�\�uɽ�*<eɽ�*<e+�n�/�Gg��	� �E�ܚ����&ꬶ�R�/���%󬷌�{�}f$W.����|̃��h�&,.�YСɽ�*<e����n��rɽ�*<eɽ�*<eɽ�*<e�����I ��(���9���wo�	h�[��w�&��^Sx=��/;~�)�D?R��9���m������VJUT���?�(<��ɽ�*<eɽ�*<eN�����K5�B���B}�k�����z�IYLy�q]�iʳ1��w�&��^Sx=��/�K��Ɛ·�z�IYLy�h���VJUT���?�(<��ɽ�*<eɽ�*<e�����^�b2�M/��J��G�I�9���g�#w�'�S 5l�[��ղ�f�!��QE���堒�c����g�#wF��@�OG�ɽ�*<eҝ[��R�ɽ�*<eɽ�*<e�r�璉�.����>W�_'����c��8;7v����ɽ�*<e�l�FD�V��jU�.2� ���c�H�hoM�Q�]�Q�Mɽ�*<e�����ɽ�*<eɽ�*<e��]/߷�W�߷G�ey�ܚ�����|�/��=1�/���%󬷌�{�}f$W.����|̃��h�&,�v�1�V�ɽ�*<e����n��rɽ�*<eɽ�*<eɽ�*<e�4ł���u}���ϖ��T�����	ɽ�*<eX��~?�W#-KB�i�`�f ��{U���g(ɽ�*<eɽ�*<eY[v�_�ɽ�*<eɽ�*<e?������|�ޒ�j\S���Γ1��#�s$����sb�F{N.J?�{�/z�E������K��(Z�ɽ�*<ex�\�uɽ�*<eɽ�*<e+�n�/�Gɕ?kV7���n�v9k���HN�E���>Է4$����sb�F{N.J��@��MQOB-�y�ɽ�*<eɽ�*<ex�\�u�~�}����7S�����F}�~RΔm����8��O6�QWk�HZ�ɽ�*<e�l�FD�V� XdJA��"C�Ӏɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<eɽ�*<e��r����<��}/���?��ɽ�*<e�Y��2�K+ҫ�0�7�/���?���h
�K=4ɽ�*<eɽ�*<eNM{9q��ɽ�*<eɽ�*<e!�T9�u�P�+H�"$-͇����i`X�F�ɽ�*<e��w�&��^<���u��D��M�N�ɽ�*<eɽ�*<e�VJUT���?�(<��ɽ�*<eɽ�*<e�]Ӟv�߷G�eyc®p"�.]��H�Q�B�/���%󬷌�{�}f��Aau�3����s�ɽ�*<eɽ�*<e����n��rɽ�*<eɽ�*<eɽ�*<e���d���xp�~�6�i�e�0ɽ�*<ea�磅"��Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���mg��gT�wQ����_���)�Ki=�Z ���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��=�wYh�ǵ��Љ�>>z�d�p�6 }m�#hL��>]�����l�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡN��Y�T��D�\å�)�}^Dz����pɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�f���y�a��b\	y`�ɽ�*<e�^1�?q�-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\U9��8P�=��O��b2�M/��J�/���%�ȣleg�׿ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc ��9t����rq��&�c���#����z:�-q26�\�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%$-͇���ג�MWz�0�\� R�E����A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%���������DC�M�T�����	ɽ�*<ea�磅"��Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���mҏ�Ba80%��;}x���ɽ�*<ei=�Z ���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��=�wYh�ǵ���c{Qb�!�Z��ɽ�*<e-&J�� ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡN��Y�T�������h���+n������pɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�f�7�D��:�M�Z��'�S 5l��^1�?q�-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\U9��8P�,{�&ZԨ�c�ޞ책�/���%��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc ��9t���\#����r�ɽ�*<esAyA/��6����[ɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%hb��e�dNl�>*�2�G���_D��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%���������DC�Mf@��S�c��.�$� ��y��5��#[���HK
ɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���m�  ƿzp��'a�y�鍕D�3�	1�$��:�Ma��͙]�ͻlU�� <�ZBg�Ҫ#MVd�ޘ ~��fɽ�*<eɽ�*<e��pJ�1
*�����{��tr��ɽ�*<eɽ�*<e^iB�j����}t�7�^*���ɽ�*<eɽ�*<e^iB�j���ڻY����L�N�����]iLɽ�*<e�%�G��>/x�kY�4V{1ɽ�*<eɽ�*<e}���5�lj��0�8�d�4V{1ɽ�*<e�/���%�`+D�o0ue'%��@�|)��t���ɽ�*<eL�@t�Z�sv/G�ˀ�ڸ�OB���c��LL�cɽ�*<eL�@t�Z�s0�{��NȈ�$r�0�2�g?�V��wɽ�*<e��U�ۄ���!���7�%����jCORuI��<ɽ�*<e�U��h���Lw��Ŝp�w���ҍ���I]ɽ�*<e7�3]N|���M��3E�c[ȈU(�ɽ�*<eɽ�*<e�.���)V�T(�<7����*���s��[ɽ�*<ed��Ję�,���,���=��Z���s��[ɽ�*<e�ߐuX�q�-�7�L���
EФ�2�H)$�e�/���%�)��;����Ј�Q�7�s-�1r����bT�>-��)ӕy0�{��NȈ��;�X���A��ͧ�>�|��
��U�ۄ����S��$�w�,\Pش��M{a����x�^6�ðU��h��f��+O���,\Pش��M{a����x�^6��7�3]N|���"�}�H�h��"'�g������
g�Z*$�V��3J�����9�����Z�l�cA�ջ�;��,�7C	d��Ję��� <�n�%W���h�J%�Y��ɽ�*<e}���5�l��p���{��%W���h�J%�Y���/���%��a'�Hs±�⳶CB���1S��M	�I�.Q"--��)ӕy0�{��NȈ�:�KD���RI��;���bT�>��U�ۄ������ �}%^Y[�\VmVW��c�=&eѼ������Xv�kɽ�*<e�/���%��8[����9(ύ��Bɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<eɽ�*<e���r�<,�����K�����]ɽ�*<e�/���%���7�1��W���[�&�E�?9D�uǎqh��gn(`m�R^0�\<efɽ�*<eɽ�*<e`ύ���#{��%B{$�`c����~�-Ȳ�N�#ɽ�*<emD�ْ�A�^_p�xqS"�3�l�\[5���d�ɽ�*<e�VJUT��� �H4%��&m(���b�{2yiglW�y���9������,(Q'�ƁQu=�U�X��~?�W#
j���?�{�/z��QT�G��J���:ɽ�*<eY[v�_�ɽ�*<eɽ�*<eA��V	{�AJ�EL�cm���fQ�΀�IPd��Qɽ�*<e�Y��2�K+)�ߙmit�`�f ��{AQ�OsJɽ�*<eɽ�*<eNM{9q��ɽ�*<eɽ�*<e!�T9�����S����]kKE��ɽ�*<eX��~?�W#
j���?�{�/z�k���C��h
�K=4ɽ�*<eY[v�_�ɽ�*<eɽ�*<e��vVK�`���;�	E\��М}��(H��u�6��/���%�Iή�%`��kC�������ʝ�u� <�t-*��h
�K=4����n��rɽ�*<eɽ�*<eɽ�*<e0��葠�Q���Д4��fMT�Ҁ����T�O�4���"#ݷIή�%`��kC����J��!㣝˻�%e�܉f��Iă�A����n��rɽ�*<eɽ�*<eɽ�*<eD���p �W"!��ٜ;���D�۳���b\	y`�ɽ�*<emD�ْ�A�^_p�x ��E��6��W��#T�.�YС�VJUT���?�(<��ɽ�*<eɽ�*<e��L��	�P�]��cR�o�O�<�ɠ)�Fɽ�*<eO��'Z
�i(�?�K��ƐΝ����%�:ɽ�*<e,4���?wɽ�*<eɽ�*<eɽ�*<e7[��İ��u}���ϖ��l�06����b��M&X��~?�W#
j���?�{�/z�k���C�w�	�6�cɽ�*<eY[v�_�ɽ�*<eɽ�*<e��vVK�`^|��]`���G�I�9��p��,ɽ�*<e[��ղ�f�}%^Y[�\Vv����W�����S�ɽ�*<eɽ�*<eҝ[��R�ɽ�*<eɽ�*<eb4�j�[���W��������h���+n�˫Y��2�K+)�ߙmit�`�f ��{�>��܎�E#L�@���ɽ�*<eNM{9q��ɽ�*<eɽ�*<e�Gy6+�$�,�IM�+�I頲wD\�w��\��ɽ�*<e�Y��2�K+)�ߙmit����
���2�h
�K=4ɽ�*<eɽ�*<eNM{9q��@82�����̟>�ĸ�����d��ve��;�d ���S3b/e�j�!I�2ɽ�*<eO��'4w��i��v[o�I�^ɽ�*<eɽ�*<e,4���?wɽ�*<eɽ�*<eɽ�*<e7[��İ��nꩠ��ʵ&�ӂ[uɽ�*<e����pɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�f#E.��#"�l��Z=�ɽ�*<e�^1�?q�-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\U9��8P�q����d��!I�2�/���%��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc ��9t�������g��h��B,k�׫�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%�)0�/ئ����#m��)/�zC�~��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%���������DC�M���,(Q'�ƁQu=�U�a�磅"��Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���mg��gT�w�W��#T�&ꬶ�Ri=�Z ���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��=�wYh�ǵ��S3b/e�j��T�O�Nd"�O��-&J�� ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡN��Y�T���R���7��$`љR�	���t�nj�'%萚 tɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�f�8��O6@��n�y֜�V��ɾ^1�?q�-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\U9��8P�G��0�@��ɽ�*<e�/���%��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc ��9t����_�av"	;��%���������ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%ז����m�b�!�Z��ɽ�*<e��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%�������~�!8��N��S���ɽ�*<e�+ �0��MK�s�Zɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���mn�W��0^�Lj}��#�˴��56i=�Z ���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��=�wYh�ǵ��nK����Mh}/Y�ɽ�*<e�����l�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡ&H'H�O�%��'X�*��U�������pɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�f#E.��#u���vQ�jɽ�*<e8\(�U�M��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\U9��8P��ܚ���ԯ�f�y��/<��\�T�h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc ��9t������(�-����)P�hx���w�E�@@ZLK|�#ɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%C�k_�pⳮ3f�d]HH��zD��}L�,4��l�ג$OJ�7��D����AP����kP�e�[�[+ɽ�*<eɽ�*<e��x��uۨ�T���]iLɽ�*<e�/���%����qBl�1nmY��
�tx�E�Bxɽ�*<e�/���%����qBl�ڸ�OB���c��LL�cɽ�*<e�/���%�6��j�.QT�'d��!3�_Fɽ�*<e�+ �0�����(T�'d��!3�_Fɽ�*<ea�+Ȳr�s�EŖڿ ˯nkB�J�tx�E�Bxɽ�*<e[a�?~��s�EŖڿ��;�X��d`���N�ɽ�*<e%"	�E׋~\�80R�|�����E_w$[��ڱ�ɽ�*<e7�3]N|���B����(c�lh��-� � x�ɽ�*<e�.���)V���-��Ǔ��x*��@M�aɽ�*<ed��Ję��j<��& �cv�A�ɽ�*<eɽ�*<e�ߐuX�q�&2}��$sN��8H��ɽ�*<e�/���%󬧁��ȉ�id=MK(�b�sN��8H��ɽ�*<e-��)ӕy0�{��NȈ|3k.sb}Hi�X&�M��aO�!�a�+Ȳr���S��$�wyu")�
B�dC�r��ɽ�*<e�U��h��|PZ��9ԁQ�onv>�v��'?�ڷI��bT�>7�3]N|� �#NS)�_Q��'�nL�n삾=Y�Aαh��T�.���)V�ֈ^��}i_Q��'�nL�n삾=Y�Aαh��Td��JęY ]}ړg��ݰI��D��L�𽼛CL��ߐuX�q�N��I-��C= 7\�&~�h����`X#Ԟ����a'�Hs�Ur���2�g�p��bxA��f���ʖ+ �0��0�{��NȈ�e�>��i�p��bxA��f���ʛ�U�ۄ����S��$�w��mf��uВ����E���bT�>�U��h���.z��7�!�қ�Bd:�6�}Zɽ�*<eY�9O=t�s��y�:3{/i�Sb�&9��̹尮l;�DhY��F�ɽ�*<e1? ��6�+t�c�K�]��s�kɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<eɽ�*<e�4����k���A�X:胮."1Do�ɽ�*<eX��~?�W#���N�^�gn(`m�R�lJ��j�<@�ͼ4���*l���űiE����nɽ�*<eɽ�*<e���Dx�v��%�6��L\�� D�(T�F(���/���%�n�>�B"�kC����I�؊nޖ�,�\�ɽ�*<e����n��ry�;Xz�����phl����?"`��%�>v;���G�I�9�[�eonD+�'V��[��ղ�fǇz��X3�v����W���D�\å�ᝄ�Dsɽ�*<eҝ[��R�ɽ�*<eɽ�*<eM�J:xc>���T�JX['����c���Gܟ�ê.ɽ�*<eyh�S
cP��ry�k��堒�c�0ڧ�AO4ɽ�*<eɽ�*<e�����ɽ�*<eɽ�*<e��]/߷�W��G�I�9mk��畬�ɽ�*<e[��ղ�fǇz��X3�v����W�"���y��ɽ�*<eɽ�*<eҝ[��R�ɽ�*<eɽ�*<em�}������u�]M���jHi��r칌,��X��~?�W#8�|q{+�?�{�/z��&�ϔ���2��Aqzɽ�*<eY[v�_�ɽ�*<eɽ�*<e��vVK�`M�L>�;>c3^Q��<8�y�P����g����!�X��~?�W#8�|q{+�?�{�/z�eg�/�b2�M/��J�h
�K=4Y[v�_�ɽ�*<eɽ�*<e�H��g澁_d�Ǹ��#��6*+�'�(.%�,aކ���jq�/���%�n�>�B"�kC�����ݮ5q.I<����<Q�]�Q�M����n��rɽ�*<eɽ�*<eɽ�*<eVd������$�!�6o�=��O����b��M&$����sb7��ɇ�F�$W.����|�z ��>�w�	�6�cɽ�*<ex�\�uɽ�*<eɽ�*<e+�n�/�G/���?����G�I�9i���!�)�49�iv ([��ղ�fǇz��X3�v����W�!&���S+�\U�>:�ɽ�*<eҝ[��R�ɽ�*<eɽ�*<em�}�����OG}Db�i���E�z�/ʛ�_�wɽ�*<e��{Y\iqS��c�Px���Y.w���`2���ɽ�*<e�VJUT���?�(<��ɽ�*<eɽ�*<e�h�z��qc�.���9r��Lj}��#�˴��56yh�S
cP��ry�k��堒�c�ɕ?kV7�'~_�~Nɽ�*<e�����ɽ�*<eɽ�*<e�t�<=��BDw��?p����`p-6�-Ȳ�N�#ɽ�*<eyh�S
cP��ry�k�\[5���d�ɽ�*<eɽ�*<eɽ�*<e�����Re|��PLz��_o�WQm$%�;���n�v9k�y�P����g�������$����sb7��ɇ�F���8��y�����ɽ�*<eɽ�*<ex�\�uɽ�*<eɽ�*<e+�n�/�G/���?���H�pf�af�w�ɽ�*<ei=�Z ���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��=�wYh�ǵ��S3b/e�jɽ�*<eɽ�*<e�����l�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡN��Y�T�!&���S+�����������pɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�fH����)x�&[�ߌ���eTq��^1�?q�-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\U9��8P�����UO`TeE+�O���0��f��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc ��9t����[�eonD+�'V�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%كY������bhF_ɽ�*<e��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%���������DC�My�P����g����!�+ �0��MK�s�Zɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���m��H�pM�L>�;>cW1	tqtV��{��Q�h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��=�wYh�ǵ��YI �_�]�ΣL%�<Y��+�2�����l�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡN��Y�T�+�T���ɽ�*<e����pɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�f�x�y�%2��Mh�]=ɽ�*<e�^1�?q�-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\U9��8P�N��S���ɽ�*<e�/���%��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc �P�~Y����z\���ɽ�*<e���z:�-q26�\�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%��(�����㗟��<�Eɽ�*<e��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%���������DC�M�/u3~�l�aކ���jqa�磅"��Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���m��G�I�9\#����r�ɽ�*<ei=�Z ���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��=�wYh�ǵ곯�	#��c�ޞ책ɽ�*<e�����E-ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡ&H'H�O�%f@��S�c��.�$� V��p�Xɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�f�8��O6Nl�>*�2�G���_DS�;��$�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\G�P�1�	��=#c?��Z�ØKϔ������!1���s�D|�����N���Q�)yū?S�$�kЈ�Q�7��b��<`�ɽ�*<e�:�<�.��0�{��NȈ�K[�k�ɽ�*<eɽ�*<eg���X���(���5V��ɽ�*<eɽ�*<eg���X0�{��NȈ��;�X��d`���N�ɽ�*<e�tO�4��S��$�w�śt�^�58���ExMɽ�*<eݵYi�f��+O���śt�^�58���ExMɽ�*<eX�&/n>�h,4���uI4M!d�>�ɽ�*<eɽ�*<e8�Cc��S��D��C��Q�onv>�v2DaZqOɽ�*<e���İ�^� = ��;��,�7C	ɽ�*<eɽ�*<ed��Ję?"(�UKx�I�tsC�0�~����~ɽ�*<e�ߐuX�q� �*�3�(�֏��ɽ�*<e�/���%󬧁��ȉ�i����7\��b�[\ɽ�*<e-��)ӕyL��P�a���ER�WV)���^Hɽ�*<e��U�ۄ���!���7�%\�j׸'��^Hɽ�*<e�U��h����R��z�F�ud�^�Ț4p�,�ɽ�*<eX�&/n>��Ҫ#MVd�e�c]���s�c�����ɽ�*<e�.���)V��ڻY����L�N��dC�r��ɽ�*<ed��Ję�#�כnp���4�MS5�w
�v.FC��ߐuX�q�3Z��Ll��np���4�MS5�w�zަ��Z�a'�Hs��9��
)��||��X���l�h��(v�cd�j�HT�[1v��zM$-����BX��hP�A~�$r�0�2K������S��$�wOhZ�ۏ�?"c���Y��ɽ�*<eݵYi����蓂s3���р�"c���Y��ɽ�*<e7�3]N|�(� ��Q'�ڑ#
�0��Bd:�6�}Zɽ�*<e�.���)V
*����䢘�9�)q���BǬ)�ɽ�*<e�8����|2w�e�Q�;��`�:�dnk�/���Z�'[P�u�ɽ�*<eɽ�*<e�
v�ƒm���X��cQ�]�Q�Mɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<eɽ�*<e^��
:�*�~�sh-�ߠwo�	h�[ɽ�*<e[��ղ�f������ܛ�*l�����R��������sk��ҝ[��R�ɽ�*<evS+ё@�˴qZ5�g�}4"{t��HN�E���>Է4X��~?�W#��	�d�?�{�/z��s��Ɩ	�q��IX;ɽ�*<ep<U˸����^1����t��.�-b|X2���H��] �, �W������˾�[(ɽ�*<e��{Y\iq���Lt�c� ��E��6�J�EL�cm�m������VJUT���?�(<��ɽ�*<eɽ�*<e�Vz�+#} �h��R�o�O�Nd"�O��ɽ�*<ex�r%=YF�����?�K��Ɛ��dsv��Zɽ�*<e,4���?wɽ�*<eɽ�*<eɽ�*<e���,hb��e�d�QWk�HZ�ɽ�*<e��{Y\iq���Lt�c�L����!��pX��ɽ�*<e�VJUT���?�(<��ɽ�*<eɽ�*<e�]Ӟv��G�I�9��rq��&�c���#�[��ղ�fǁ����=�v����W���R���7���՞WS�ɽ�*<eҝ[��R�ɽ�*<eɽ�*<e��{P���� <�t-*���G�I�9/���?��..+`��[��ղ�fǁ����=�v����W���P�6;7}��]oT5��ɽ�*<eҝ[��R�ɽ�*<eɽ�*<e���U�&4��%e�܉��+ά���������J�\� R�E��X��~?�W#��	�d�?�{�/z�wM�.�����$�c>y�Dɽ�*<eY[v�_�ɽ�*<eɽ�*<eA��V	{�A�W��#T���0�7��P�6;7}49�iv (�Y��2�K+�I�\�m��`�f ��{�f>;�݃�\U�>:�ɽ�*<eNM{9q��ɽ�*<eɽ�*<e!�T9�u�P�+H�"hb��e�dB�$Dɽ�*<e��{Y\iq���Lt�c�L����^|��]`��h
�K=4�VJUT���?�(<��ɽ�*<eɽ�*<e�]Ӟv�߷G�ey&6��u48ɽ�*<e�/���%�|2w�e�Q��kC����̾���ܔ7]��s�kɽ�*<e����n��rɽ�*<eɽ�*<eɽ�*<eU�Z�H� �-�!Ɖc�㗟��<�Eɽ�*<ex�r%=YF�����?�ч�t}�,�IM�+�IQOB-�y�,4���?wɽ�*<eɽ�*<eɽ�*<e�|.���s��@B�#h��4�(T�F(��ɽ�*<ex�r%=YF��k�UhU�Gޖ�,�\�ɽ�*<eɽ�*<e,4���?wMͿ���q�����&�R@I�K�E���D�M�N�頲wD\�/���?��ɽ�*<e�Y��2�K+�I�\�m�ʿ�P�6;7}�&ZReX�ɽ�*<eɽ�*<eNM{9q��ɽ�*<eɽ�*<e!�T9�u�P�+H�"$-͇���ה'd����ɽ�*<e��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%���������DC�Mi�e�0ɽ�*<ea�磅"��Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���m��H�p^|��]`�ɽ�*<ei=�Z ���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��=�wYh�ǵ��Љ�>>z�c��<��iP��[P�����l�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡN��Y�T��A������s �� rA�Uc�_:ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�f9+v�r�ô�˾�[(ɽ�*<e�^1�?q�-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\U9��8P�V�3yn�3y֜�V����/���%��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc ��9t���/���?��..+`�����z:�-q26�\�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%[������ <�t-*�ɽ�*<e(�B)�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%���������DC�M*����>�W��#T�aD���^�aQ�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���m�)��H�6��D�j�)Iɽ�*<ei=�Z ���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��=�wYh�ǵ�+��,�]�D��~��ɽ�*<e�����l�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡN��Y�T�z\���ɽ�*<e����pɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�f܁:ze��d��;}x���ɽ�*<eS�;��$�Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\U9��8P�S���Γ1��#�s�/���%��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc ��9t���_tp�n�.]\� R�E�ի�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%B}�k���u���vQ�jɽ�*<e��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%���������DC�M��'X�*��U����:�<�.�ؙCB"��,#ɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���m��G�I�9���(�-����)P�hx�E���G�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��=�wYh�ǵ��YI �_��f�y������&8_K��c��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡ����Ve:�X��\��ݑ��/�^�L�Lr)��ש0��b=��K�X}(�K�r�UP����yu")�
B����]iLɽ�*<e�i��K���.z��7��1�p%�F�ɽ�*<eɽ�*<e-&�
:lݲf��+O��P�.a7)�ɽ�*<eɽ�*<e-&�
:lݲ|PZ��9ԁQ�onv>�v2DaZqOɽ�*<e�
���Wϓ��g��b��<�Z�%�tx�E�Bxɽ�*<eB�j�^9TŤ�м�U�<�Z�%�tx�E�Bxɽ�*<e�dtD<]�<�y5c@����&�Ī;��ɽ�*<eɽ�*<e�A����׏��w��C����L�N�����]iLɽ�*<e�%����F_hHbJ�3��x�K��ɽ�*<e�/���%󬧁��ȉ�iLD�d��9__n�X�t�ɽ�*<e-��)ӕyL��P�a�����>Sp�ޞx�-�ɽ�*<e��U�ۄ���!���7�%#N7Q���N�dh1zɽ�*<e�U��h���Lw�羈�g���.�Dz�.�ɽ�*<e7�3]N|��r)d`b��\�()�Ľ.�Dz�.�ɽ�*<e�.���)Vi}^�k�fU���Ɔ[7����ɽ�*<e�dtD<]�<�AP����k ��y$���>�|��
ɽ�*<e�ߐuX�q�ڸ�OB��ur�$��s�c������/���%��a'�Hs���`�^+�>�JƬӣ�a
k��K1<NSmr�c���(��`�^+�>�JƬӣ�a
k��K1��-�y�Y���S��$�w��}hm�As�FJ������ (�ҬR�n�f���M���Y^�+������V,�U��|�����E_��Ύ���"�}�H�h\rһ�ޏJ=P�P9Qɽ�*<eB�j�^9
QX������<����J=P�P9Qɽ�*<ed��Ję���Ϧt�*NZ�g�BǬ)�ɽ�*<e�ߐuX�q��uۨ�T�s�g��8Z	�I�.Q"-�/���%󬱖����(��Jnj��IK�vv��O�ơ���a'ѳ��w��ɽ�*<eɽ�*<e��=!��(2��p�ɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<��ɽ�*<e:j���+�oaf�	��,��/�=X]ɽ�*<eɽ�*<emD�ْ�dh89QN��hz�;3��PY���F��
�W���[�&���2�%?�(<��ɽ�*<e��_��l���<I}���G�I�9w��\��ɽ�*<e[��ղ�f�ڇ��C�v����W����
���2�h
�K=4ɽ�*<eVӥRysL_ �1J�`���u@�:4j�ק�	��� 4���:o�W��JW����sp��/���%�;K�Raz�kC�����o�2��vc6%8�s���Q�]�Q�M����n��rɽ�*<eɽ�*<eɽ�*<e��"�m҂B�1ci��)�<�;ɽ�*<e$����sbt���̌$W.����|�z ��>��h
�K=4ɽ�*<ex�\�uɽ�*<eɽ�*<e+�n�/�Gg��	� �E�ܚ����&ꬶ�R�/���%�;K�Raz�kC�����z��=S�w��Rdɽ�*<e����n��rɽ�*<eɽ�*<eɽ�*<e�����I ��(���9���wo�	h�[��{Y\iq��;�TL����M�L>�;>cc��R��Mb�VJUT���?�(<��ɽ�*<eɽ�*<eN�����K5�B���B}�k�����z�IYLy�q]�iʳ1��{Y\iq��;�T2� ���_d�Ǹ��..
A����VJUT���?�(<��ɽ�*<eɽ�*<e�����^�b2�M/��J��G�I�9���g�#w�'�S 5l�[��ղ�f�ڇ��C�v����W��Д�٪,EWP���ɽ�*<eҝ[��R�ɽ�*<eɽ�*<e�r�璉�.����>W�_'����c��8;7v����ɽ�*<eyh�S
cP�Ɖ�D��0L�堒�c�/���?���h
�K=4ɽ�*<e�����ɽ�*<eɽ�*<e��]/߷�W�߷G�ey�ܚ�����|�/��=1�/���%�;K�Raz�kC�����z��=D��M�N�ɽ�*<e����n��rɽ�*<eɽ�*<eɽ�*<e�4ł���u}���ϖ��T�����	ɽ�*<eX��~?�W#��Jnj��?�{�/z����c��kQ�]�Q�Mɽ�*<eY[v�_�ɽ�*<eɽ�*<e?������|�ޒ�j\S���Γ1��#�s$����sbt���̌$W.����|�� �"y&�sn5&;�Q�]�Q�Mx�\�uɽ�*<eɽ�*<e+�n�/�Gɕ?kV7���n�v9k���HN�E���>Է4$����sbt���̌/���>;�#	�q��IX;ɽ�*<eɽ�*<ex�\�u�~�}����7S�����F}�~RΔm���#E.��#5�'��,��ɽ�*<eyh�S
cP�{�p���c�H�hoM�Q�]�Q�Mɽ�*<eɽ�*<e�����ɽ�*<eɽ�*<e��]/߷�W�߷G�eyq����d�ɽ�*<e�/���%��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc ��9t���"�d�;�ɽ�*<e������ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%$-͇����i`X�F�ɽ�*<e��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%���������DC�Mz`��'9�)/�zC�~a�磅"��Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���mg��gT�w<u��rnN�-����ngMܵ�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��=�wYh�ǵ�I��u+��(W����sp�ɽ�*<e�����l�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡN��Y�T�Д�٪,<Y��+�2����pɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�f#E.��#��z�IYLy�q]�iʳ1S�;��$�Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\U9��8P�ZQ�R�"=�5�7��dh�/���%�ȣleg�׿ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc ��9t���;����L��bhF_������ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%du���1�DhY��F�ɽ�*<e��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%���������DC�M��0ך��0��F��X�a�磅"��Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���mҏ�Ba80%��;}x���ɽ�*<ei=�Z ���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��=�wYh�ǵ���c{Qb�!�Z��ɽ�*<e-&J�� ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡN��Y�T�������h���+n������pɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�f�7�D��:�M�Z��'�S 5l��^1�?q�-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\U9��8P�,{�&ZԨ�c�ޞ책�/���%��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc ��9t���\#����r�ɽ�*<esAyA/��6����[ɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%hb��e�dNl�>*�2�G���_D��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%���������DC�Mf@��S�c��.�$� ��y��5��#[���HK
ɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���m�  ƿzp��'a�y�鍕D�3�	1�$��:�Ma��͙]�ͻlU�� <�ZBg�Ҫ#MVd�ޘ ~��fɽ�*<eɽ�*<e��pJ�1
*�����{��tr��ɽ�*<eɽ�*<e^iB�j����}t�7�^*���ɽ�*<eɽ�*<e^iB�j���ڻY����L�N�����]iLɽ�*<e�%�G��>/x�kY�4V{1ɽ�*<eɽ�*<e}���5�lj��0�8�d�4V{1ɽ�*<e�/���%�`+D�o0ue'%��@�|)��t���ɽ�*<eL�@t�Z�sv/G�ˀ�ڸ�OB���c��LL�cɽ�*<eL�@t�Z�s0�{��NȈ�$r�0�2�g?�V��wɽ�*<e��U�ۄ���!���7�%����jCORuI��<ɽ�*<e�U��h���Lw��Ŝp�w���ҍ���I]ɽ�*<e7�3]N|���M��3E�c[ȈU(�ɽ�*<eɽ�*<e�.���)V�T(�<7����*���s��[ɽ�*<ed��Ję�,���,���=��Z���s��[ɽ�*<e�ߐuX�q�-�7�L���
EФ�2�H)$�e�/���%�)��;����Ј�Q�7�s-�1r����bT�>-��)ӕy0�{��NȈ��;�X���A��ͧ�>�|��
��U�ۄ����S��$�w�,\Pش��M{a����x�^6�ðU��h��f��+O���,\Pش��M{a����x�^6��7�3]N|���"�}�H�h��"'�g������
g�Z*$�V��3J�����9�����Z�l�cA�ջ�;��,�7C	d��Ję��� <�n�%W���h�J%�Y��ɽ�*<e}���5�l��p���{��%W���h�J%�Y���/���%��a'�Hs±�⳶CB���1S��M	�I�.Q"--��)ӕy0�{��NȈ�:�KD���RI��;���bT�>��U�ۄ������ �������mVW��c�=&eѼ������Xv�kɽ�*<e�/���%��8[����9(ύ��Bɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<eɽ�*<e���r�<,�����K�����]ɽ�*<e�/���%���7�1��W���[�&�E�?9D�uǎqh��gn(`m�R^0�\<efɽ�*<eɽ�*<e`ύ���#{��%B{$�`c����~�-Ȳ�N�#ɽ�*<e��{Y\iq��Ժ��h�qS"�3�l�\[5���d�ɽ�*<e�VJUT��� �H4%��&m(���b�{2yiglW�y���9������,(Q'�ƁQu=�U�X��~?�W#|m9T�g�R?�{�/z��QT�G��J���:ɽ�*<eY[v�_�ɽ�*<eɽ�*<eA��V	{�AJ�EL�cm���fQ�΀�IPd��Qɽ�*<e�Y��2�K+���]-��`�f ��{AQ�OsJɽ�*<eɽ�*<eNM{9q��ɽ�*<eɽ�*<e!�T9�����S����]kKE��ɽ�*<eX��~?�W#|m9T�g�R?�{�/z�k���C��h
�K=4ɽ�*<eY[v�_�ɽ�*<eɽ�*<e��vVK�`���;�	E\��М}��(H��u�6��/���%󬖸3����kC�������ʝ�u� <�t-*��h
�K=4����n��rɽ�*<eɽ�*<eɽ�*<e0��葠�Q���Д4��fMT�Ҁ����T�O�4���"#ݷ��3����kC����J��!㣝˻�%e�܉f��Iă�A����n��rɽ�*<eɽ�*<eɽ�*<eD���p �W"!��ٜ;���D�۳���b\	y`�ɽ�*<e��{Y\iq��Ժ��h� ��E��6��W��#T�.�YС�VJUT���?�(<��ɽ�*<eɽ�*<e��L��	�P�]��cR�o�O�<�ɠ)�Fɽ�*<ex�r%=YF�N'������K��ƐΝ����%�:ɽ�*<e,4���?wɽ�*<eɽ�*<eɽ�*<e7[��İ��u}���ϖ��l�06����b��M&X��~?�W#|m9T�g�R?�{�/z�k���C�w�	�6�cɽ�*<eY[v�_�ɽ�*<eɽ�*<e��vVK�`^|��]`���G�I�9��p��,ɽ�*<e[��ղ�f�������v����W�����S�ɽ�*<eɽ�*<eҝ[��R�ɽ�*<eɽ�*<eb4�j�[���W��������h���+n�˫Y��2�K+���]-��`�f ��{�>��܎�E#L�@���ɽ�*<eNM{9q��ɽ�*<eɽ�*<e�Gy6+�$�,�IM�+�I頲wD\�w��\��ɽ�*<e�Y��2�K+���]-�����
���2�h
�K=4ɽ�*<eɽ�*<eNM{9q��@82�����̟>�ĸ�����d��ve��;�d ���S3b/e�j�!I�2ɽ�*<ex�r%=YF�m5�C��e�v[o�I�^ɽ�*<eɽ�*<e,4���?wɽ�*<eɽ�*<eɽ�*<e7[��İ��nꩠ��ʵ&�ӂ[uɽ�*<e����pɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�f#E.��#"�l��Z=�ɽ�*<e�^1�?q�-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\U9��8P�q����d��!I�2�/���%��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc ��9t�������g��h��B,k�׫�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%�)0�/ئ����#m��)/�zC�~��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%���������DC�M���,(Q'�ƁQu=�U�a�磅"��Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���mg��gT�w�W��#T�&ꬶ�Ri=�Z ���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��=�wYh�ǵ��S3b/e�j��T�O�Nd"�O��-&J�� ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡN��Y�T���R���7��$`љR�	���t�nj�'%萚 tɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�f�8��O6@��n�y֜�V��ɾ^1�?q�-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\U9��8P�G��0�@��ɽ�*<e�/���%��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc ��9t����_�av"	;��%���������ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%ז����m�b�!�Z��ɽ�*<e��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%�������~�!8��N��S���ɽ�*<e�+ �0��MK�s�Zɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���mn�W��0^�Lj}��#�˴��56i=�Z ���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��=�wYh�ǵ��nK����Mh}/Y�ɽ�*<e�����l�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡ&H'H�O�%��'X�*��U�������pɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�f#E.��#u���vQ�jɽ�*<e8\(�U�M��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\U9��8P��ܚ���ԯ�f�y��/<��\�T�h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc ��9t������(�-����)P�hx���w�E�@@ZLK|�#ɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%C�k_�pⳮ3f�d]HH��zD��}L�,4��l�ג$OJ�7��D����AP����kP�e�[�[+ɽ�*<eɽ�*<e��x��uۨ�T���]iLɽ�*<e�/���%����qBl�1nmY��
�tx�E�Bxɽ�*<e�/���%����qBl�ڸ�OB���c��LL�cɽ�*<e�/���%�6��j�.QT�'d��!3�_Fɽ�*<e�+ �0�����(T�'d��!3�_Fɽ�*<ea�+Ȳr�s�EŖڿ ˯nkB�J�tx�E�Bxɽ�*<e[a�?~��s�EŖڿ��;�X��d`���N�ɽ�*<e%"	�E׋~\�80R�|�����E_w$[��ڱ�ɽ�*<e7�3]N|���B����(c�lh��-� � x�ɽ�*<e�.���)V���-��Ǔ��x*��@M�aɽ�*<ed��Ję��j<��& �cv�A�ɽ�*<eɽ�*<e�ߐuX�q�&2}��$sN��8H��ɽ�*<e�/���%󬧁��ȉ�id=MK(�b�sN��8H��ɽ�*<e-��)ӕy0�{��NȈ|3k.sb}Hi�X&�M��aO�!�a�+Ȳr���S��$�wyu")�
B�dC�r��ɽ�*<e�U��h��|PZ��9ԁQ�onv>�v��'?�ڷI��bT�>7�3]N|� �#NS)�_Q��'�nL�n삾=Y�Aαh��T�.���)V�ֈ^��}i_Q��'�nL�n삾=Y�Aαh��Td��JęY ]}ړg��ݰI��D��L�𽼛CL��ߐuX�q�N��I-��C= 7\�&~�h����`X#Ԟ����a'�Hs�Ur���2�g�p��bxA��f���ʖ+ �0��0�{��NȈ�e�>��i�p��bxA��f���ʛ�U�ۄ����S��$�w��mf��uВ����E���bT�>�U��h���.z��7�!�қ�Bd:�6�}Zɽ�*<eY�9O=t�s��y��l�,�`��Sb�&9��̹尮l;�DhY��F�ɽ�*<e1? ��6�+t�c�K�]��s�kɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<eɽ�*<e�4����k���A�X:胮."1Do�ɽ�*<eX��~?�W#���N�^�gn(`m�R�lJ��j�<@�ͼ4���*l���űiE����nɽ�*<eɽ�*<e���Dx�v��%�6��L\�� D�(T�F(���/���%���f�|L�kC����I�؊nޖ�,�\�ɽ�*<e����n��ry�;Xz�����phl����?"`��%�>v;���G�I�9�[�eonD+�'V��[��ղ�fǕpᓖC�v����W���D�\å�ᝄ�Dsɽ�*<eҝ[��R�ɽ�*<eɽ�*<eM�J:xc>���T�JX['����c���Gܟ�ê.ɽ�*<eyh�S
cP�����N�B�堒�c�0ڧ�AO4ɽ�*<eɽ�*<e�����ɽ�*<eɽ�*<e��]/߷�W��G�I�9mk��畬�ɽ�*<e[��ղ�fǕpᓖC�v����W�"���y��ɽ�*<eɽ�*<eҝ[��R�ɽ�*<eɽ�*<em�}������u�]M���jHi��r칌,��X��~?�W#;i���`C>?�{�/z��&�ϔ���2��Aqzɽ�*<eY[v�_�ɽ�*<eɽ�*<e��vVK�`M�L>�;>c3^Q��<8�y�P����g����!�X��~?�W#;i���`C>?�{�/z�eg�/�b2�M/��J�h
�K=4Y[v�_�ɽ�*<eɽ�*<e�H��g澁_d�Ǹ��#��6*+�'�(.%�,aކ���jq�/���%���f�|L�kC�����ݮ5q.I<����<Q�]�Q�M����n��rɽ�*<eɽ�*<eɽ�*<eVd������$�!�6o�=��O����b��M&$����sb(�2Y�ǫ$W.����|�z ��>�w�	�6�cɽ�*<ex�\�uɽ�*<eɽ�*<e+�n�/�G/���?����G�I�9i���!�)�49�iv ([��ղ�fǕpᓖC�v����W�!&���S+�\U�>:�ɽ�*<eҝ[��R�ɽ�*<eɽ�*<em�}�����OG}Db�i���E�z�/ʛ�_�wɽ�*<e��{Y\iqd������x���Y.w���`2���ɽ�*<e�VJUT���?�(<��ɽ�*<eɽ�*<e�h�z��qc�.���9r��Lj}��#�˴��56yh�S
cP�����N�B�堒�c�ɕ?kV7�'~_�~Nɽ�*<e�����ɽ�*<eɽ�*<e�t�<=��BDw��?p����`p-6�-Ȳ�N�#ɽ�*<eyh�S
cP�����N�B\[5���d�ɽ�*<eɽ�*<eɽ�*<e�����Re|��PLz��_o�WQm$%�;���n�v9k�y�P����g�������$����sb(�2Y�ǫ��8��y�����ɽ�*<eɽ�*<ex�\�uɽ�*<eɽ�*<e+�n�/�G/���?���H�pf�af�w�ɽ�*<ei=�Z ���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��=�wYh�ǵ��S3b/e�jɽ�*<eɽ�*<e�����l�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡN��Y�T�!&���S+�����������pɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�fH����)x�&[�ߌ���eTq��^1�?q�-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\U9��8P�����UO`TeE+�O���0��f��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc ��9t����[�eonD+�'V�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%كY������bhF_ɽ�*<e��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%���������DC�My�P����g����!�+ �0��MK�s�Zɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���m��H�pM�L>�;>cW1	tqtV��{��Q�h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��=�wYh�ǵ��YI �_�]�ΣL%�<Y��+�2�����l�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡN��Y�T�+�T���ɽ�*<e����pɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�f�x�y�%2��Mh�]=ɽ�*<e�^1�?q�-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\U9��8P�N��S���ɽ�*<e�/���%��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc �P�~Y����z\���ɽ�*<e���z:�-q26�\�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%��(�����㗟��<�Eɽ�*<e��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%���������DC�M�/u3~�l�aކ���jqa�磅"��Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���m��G�I�9\#����r�ɽ�*<ei=�Z ���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��=�wYh�ǵ곯�	#��c�ޞ책ɽ�*<e�����E-ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡ&H'H�O�%f@��S�c��.�$� V��p�Xɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�f�8��O6Nl�>*�2�G���_DS�;��$�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\G�P�1�	��=#c?��Z�ØKϔ������!1���s�D|�����N���Q�)yū?S�$�kЈ�Q�7��b��<`�ɽ�*<e�:�<�.��0�{��NȈ�K[�k�ɽ�*<eɽ�*<eg���X���(���5V��ɽ�*<eɽ�*<eg���X0�{��NȈ��;�X��d`���N�ɽ�*<e�tO�4��S��$�w�śt�^�58���ExMɽ�*<eݵYi�f��+O���śt�^�58���ExMɽ�*<eX�&/n>�h,4���uI4M!d�>�ɽ�*<eɽ�*<e8�Cc��S��D��C��Q�onv>�v2DaZqOɽ�*<e���İ�^� = ��;��,�7C	ɽ�*<eɽ�*<ed��Ję?"(�UKx�I�tsC�0�~����~ɽ�*<e�ߐuX�q� �*�3�(�֏��ɽ�*<e�/���%󬧁��ȉ�i����7\��b�[\ɽ�*<e-��)ӕyL��P�a���ER�WV)���^Hɽ�*<e��U�ۄ���!���7�%\�j׸'��^Hɽ�*<e�U��h����R��z�F�ud�^�Ț4p�,�ɽ�*<eX�&/n>��Ҫ#MVd�e�c]���s�c�����ɽ�*<e�.���)V��ڻY����L�N��dC�r��ɽ�*<ed��Ję�#�כnp���4�MS5�w
�v.FC��ߐuX�q�3Z��Ll��np���4�MS5�w�zަ��Z�a'�Hs��9��
)��||��X���l�h��(v�cd�j�HT�[1v��zM$-����BX��hP�A~�$r�0�2K������S��$�wOhZ�ۏ�?"c���Y��ɽ�*<eݵYi����蓂s3���р�"c���Y��ɽ�*<e7�3]N|�(� ��Q'�ڑ#
�0��Bd:�6�}Zɽ�*<e�.���)V
*����䢘�9�)q���BǬ)�ɽ�*<e�8�����/�ӄi�4;��`�:�dnk�/���Z�'[P�u�ɽ�*<eɽ�*<e�
v�ƒm���X��cQ�]�Q�Mɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<eɽ�*<e^��
:�*�~�sh-�ߠwo�	h�[ɽ�*<e[��ղ�f������ܛ�*l�����R��������sk��ҝ[��R�ɽ�*<evS+ё@�˴qZ5�g�}4"{t��HN�E���>Է4X��~?�W#e���I?�{�/z��s��Ɩ	�q��IX;ɽ�*<ep<U˸����^1����t��.�-b|X2���H��] �, �W������˾�[(ɽ�*<e��{Y\iq�f�� ��E��6�J�EL�cm�m������VJUT���?�(<��ɽ�*<eɽ�*<e�Vz�+#} �h��R�o�O�Nd"�O��ɽ�*<ex�r%=YF�2h�L�&�_�K��Ɛ��dsv��Zɽ�*<e,4���?wɽ�*<eɽ�*<eɽ�*<e���,hb��e�d�QWk�HZ�ɽ�*<e��{Y\iq�f��L����!��pX��ɽ�*<e�VJUT���?�(<��ɽ�*<eɽ�*<e�]Ӟv��G�I�9��rq��&�c���#�[��ղ�f�H���5�v����W���R���7���՞WS�ɽ�*<eҝ[��R�ɽ�*<eɽ�*<e��{P���� <�t-*���G�I�9/���?��..+`��[��ղ�f�H���5�v����W���P�6;7}��]oT5��ɽ�*<eҝ[��R�ɽ�*<eɽ�*<e���U�&4��%e�܉��+ά���������J�\� R�E��X��~?�W#e���I?�{�/z�wM�.�����$�c>y�Dɽ�*<eY[v�_�ɽ�*<eɽ�*<eA��V	{�A�W��#T���0�7��P�6;7}49�iv (�Y��2�K+I�b�H�`�f ��{�f>;�݃�\U�>:�ɽ�*<eNM{9q��ɽ�*<eɽ�*<e!�T9�u�P�+H�"hb��e�dB�$Dɽ�*<e��{Y\iq�f��L����^|��]`��h
�K=4�VJUT���?�(<��ɽ�*<eɽ�*<e�]Ӟv�߷G�ey&6��u48ɽ�*<e�/���%��/�ӄi�4�kC����̾���ܔ7]��s�kɽ�*<e����n��rɽ�*<eɽ�*<eɽ�*<eU�Z�H� �-�!Ɖc�㗟��<�Eɽ�*<ex�r%=YF�2h�L�&�_�ч�t}�,�IM�+�IQOB-�y�,4���?wɽ�*<eɽ�*<eɽ�*<e�|.���s��@B�#h��4�(T�F(��ɽ�*<ex�r%=YF���q�6x�ޖ�,�\�ɽ�*<eɽ�*<e,4���?wMͿ���q�����&�R@I�K�E���D�M�N�頲wD\�/���?��ɽ�*<e�Y��2�K+I�b�H濘P�6;7}�&ZReX�ɽ�*<eɽ�*<eNM{9q��ɽ�*<eɽ�*<e!�T9�u�P�+H�"$-͇���ה'd����ɽ�*<e��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%���������DC�Mi�e�0ɽ�*<ea�磅"��Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���m��H�p^|��]`�ɽ�*<ei=�Z ���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��=�wYh�ǵ��Љ�>>z�c��<��iP��[P�����l�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡN��Y�T��A������s �� rA�Uc�_:ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�f9+v�r�ô�˾�[(ɽ�*<e�^1�?q�-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\U9��8P�V�3yn�3y֜�V����/���%��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc ��9t���/���?��..+`�����z:�-q26�\�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%[������ <�t-*�ɽ�*<e(�B)�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%���������DC�M*����>�W��#T�aD���^�aQ�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���m�)��H�6��D�j�)Iɽ�*<ei=�Z ���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��=�wYh�ǵ�+��,�]�D��~��ɽ�*<e�����l�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡN��Y�T�z\���ɽ�*<e����pɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�f܁:ze��d��;}x���ɽ�*<eS�;��$�Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\U9��8P�S���Γ1��#�s�/���%��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc ��9t���_tp�n�.]\� R�E�ի�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%B}�k���u���vQ�jɽ�*<e��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%���������DC�M��'X�*��U����:�<�.�ؙCB"��,#ɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���m��G�I�9���(�-����)P�hx�E���G�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��=�wYh�ǵ��YI �_��f�y������&8_K��c��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡ����Ve:�X��\��ݑ��/�^�L�Lr)��ש0��b=��K�X}(�K�r�UP����yu")�
B����]iLɽ�*<e�i��K���.z��7��1�p%�F�ɽ�*<eɽ�*<e-&�
:lݲf��+O��P�.a7)�ɽ�*<eɽ�*<e-&�
:lݲ|PZ��9ԁQ�onv>�v2DaZqOɽ�*<e�
���Wϓ��g��b��<�Z�%�tx�E�Bxɽ�*<eB�j�^9TŤ�м�U�<�Z�%�tx�E�Bxɽ�*<e�dtD<]�<�y5c@����&�Ī;��ɽ�*<eɽ�*<e�A����׏��w��C����L�N�����]iLɽ�*<e�%����F_hHbJ�3��x�K��ɽ�*<e�/���%󬧁��ȉ�iLD�d��9__n�X�t�ɽ�*<e-��)ӕyL��P�a�����>Sp�ޞx�-�ɽ�*<e��U�ۄ���!���7�%#N7Q���N�dh1zɽ�*<e�U��h���Lw�羈�g���.�Dz�.�ɽ�*<e7�3]N|��r)d`b��\�()�Ľ.�Dz�.�ɽ�*<e�.���)Vi}^�k�fU���Ɔ[7����ɽ�*<e�dtD<]�<�AP����k ��y$���>�|��
ɽ�*<e�ߐuX�q�ڸ�OB��ur�$��s�c������/���%��a'�Hs���`�^+�>�JƬӣ�a
k��K1<NSmr�c���(��`�^+�>�JƬӣ�a
k��K1��-�y�Y���S��$�w��}hm�As�FJ������ (�ҬR�n�f���M���Y^�+������V,�U��|�����E_��Ύ���"�}�H�h\rһ�ޏJ=P�P9Qɽ�*<eB�j�^9
QX������<����J=P�P9Qɽ�*<ed��Ję���Ϧt�*NZ�g�BǬ)�ɽ�*<e�ߐuX�q��uۨ�T�s�g��8Z	�I�.Q"-�/���%󬱖����(�`���$��IK�vv��O�ơ���a'ѳ��w��ɽ�*<eɽ�*<e��=!��(2��p�ɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<��ɽ�*<e:j���+�oaf�	��,��/�=X]ɽ�*<eɽ�*<emD�ْ�dh89QN��hz�;3��PY���F��
�W���[�&���2�%?�(<��ɽ�*<e��_��l���<I}���G�I�9w��\��ɽ�*<e[��ղ�f��\�m0a�v����W����
���2�h
�K=4ɽ�*<eVӥRysL_ �1J�`���u@�:4j�ק�	��� 4���:o�W��JW����sp��/���%���?��B��kC�����o�2��vc6%8�s���Q�]�Q�M����n��rɽ�*<eɽ�*<eɽ�*<e��"�m҂B�1ci��)�<�;ɽ�*<e$����sb�s7�}��$W.����|�z ��>��h
�K=4ɽ�*<ex�\�uɽ�*<eɽ�*<e+�n�/�Gg��	� �E�ܚ����&ꬶ�R�/���%���?��B��kC�����z��=S�w��Rdɽ�*<e����n��rɽ�*<eɽ�*<eɽ�*<e�����I ��(���9���wo�	h�[��{Y\iq*��ř%(L����M�L>�;>cc��R��Mb�VJUT���?�(<��ɽ�*<eɽ�*<eN�����K5�B���B}�k�����z�IYLy�q]�iʳ1��{Y\iq*��ř%(2� ���_d�Ǹ��..
A����VJUT���?�(<��ɽ�*<eɽ�*<e�����^�b2�M/��J��G�I�9���g�#w�'�S 5l�[��ղ�f��\�m0a�v����W��Д�٪,EWP���ɽ�*<eҝ[��R�ɽ�*<eɽ�*<e�r�璉�.����>W�_'����c��8;7v����ɽ�*<eyh�S
cP�r)1�ڹ��堒�c�/���?���h
�K=4ɽ�*<e�����ɽ�*<eɽ�*<e��]/߷�W�߷G�ey�ܚ�����|�/��=1�/���%���?��B��kC�����z��=D��M�N�ɽ�*<e����n��rɽ�*<eɽ�*<eɽ�*<e�4ł���u}���ϖ��T�����	ɽ�*<eX��~?�W#�`���$��?�{�/z����c��kQ�]�Q�Mɽ�*<eY[v�_�ɽ�*<eɽ�*<e?������|�ޒ�j\S���Γ1��#�s$����sb�s7�}��$W.����|�� �"y&�sn5&;�Q�]�Q�Mx�\�uɽ�*<eɽ�*<e+�n�/�Gɕ?kV7���n�v9k���HN�E���>Է4$����sb�s7�}��/���>;�#	�q��IX;ɽ�*<eɽ�*<ex�\�u�~�}����7S�����F}�~RΔm���#E.��#5�'��,��ɽ�*<eyh�S
cP��tw
�Z�c�H�hoM�Q�]�Q�Mɽ�*<eɽ�*<e�����ɽ�*<eɽ�*<e��]/߷�W�߷G�eyq����d�ɽ�*<e�/���%��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc ��9t���"�d�;�ɽ�*<e������ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%$-͇����i`X�F�ɽ�*<e��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%���������DC�Mz`��'9�)/�zC�~a�磅"��Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���mg��gT�w<u��rnN�-����ngMܵ�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��=�wYh�ǵ�I��u+��(W����sp�ɽ�*<e�����l�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡN��Y�T�Д�٪,<Y��+�2����pɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�f#E.��#��z�IYLy�q]�iʳ1S�;��$�Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\U9��8P�ZQ�R�"=�5�7��dh�/���%�ȣleg�׿ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc ��9t���;����L��bhF_������ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%du���1�DhY��F�ɽ�*<e��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%���������DC�M��0ך��0��F��X�a�磅"��Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���mҏ�Ba80%��;}x���ɽ�*<ei=�Z ���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��=�wYh�ǵ���c{Qb�!�Z��ɽ�*<e-&J�� ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡN��Y�T�������h���+n������pɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�f�7�D��:�M�Z��'�S 5l��^1�?q�-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\U9��8P�,{�&ZԨ�c�ޞ책�/���%��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc ��9t���\#����r�ɽ�*<esAyA/��6����[ɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%hb��e�dNl�>*�2�G���_D��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%���������DC�Mf@��S�c��.�$� ��y��5��#[���HK
ɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���m�  ƿzp��'a�y�鍕D�3�	1�$��:�Ma��͙]�ͻlU�� <�ZBg�Ҫ#MVd�ޘ ~��fɽ�*<eɽ�*<e��pJ�1
*�����{��tr��ɽ�*<eɽ�*<e^iB�j����}t�7�^*���ɽ�*<eɽ�*<e^iB�j���ڻY����L�N�����]iLɽ�*<e�%�G��>/x�kY�4V{1ɽ�*<eɽ�*<e}���5�lj��0�8�d�4V{1ɽ�*<e�/���%�`+D�o0ue'%��@�|)��t���ɽ�*<eL�@t�Z�sv/G�ˀ�ڸ�OB���c��LL�cɽ�*<eL�@t�Z�s0�{��NȈ�$r�0�2�g?�V��wɽ�*<e��U�ۄ���!���7�%����jCORuI��<ɽ�*<e�U��h���Lw��Ŝp�w���ҍ���I]ɽ�*<e7�3]N|���M��3E�c[ȈU(�ɽ�*<eɽ�*<e�.���)V�T(�<7����*���s��[ɽ�*<ed��Ję�,���,���=��Z���s��[ɽ�*<e�ߐuX�q�-�7�L���
EФ�2�H)$�e�/���%�)��;����Ј�Q�7�s-�1r����bT�>-��)ӕy0�{��NȈ��;�X���A��ͧ�>�|��
��U�ۄ����S��$�w�,\Pش��M{a����x�^6�ðU��h��f��+O���,\Pش��M{a����x�^6��7�3]N|���"�}�H�h��"'�g������
g�Z*$�V��3J�����9�����Z�l�cA�ջ�;��,�7C	d��Ję��� <�n�%W���h�J%�Y��ɽ�*<e}���5�l��p���{��%W���h�J%�Y���/���%��a'�Hs±�⳶CB���1S��M	�I�.Q"--��)ӕy0�{��NȈ�:�KD���RI��;���bT�>��U�ۄ������ � �D�O�h>mVW��c�=&eѼ������Xv�kɽ�*<e�/���%��8[����9(ύ��Bɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<eɽ�*<e���r�<,�����K�����]ɽ�*<e�/���%���7�1��W���[�&�E�?9D�uǎqh��gn(`m�R^0�\<efɽ�*<eɽ�*<e`ύ���#{��%B{$�`c����~�-Ȳ�N�#ɽ�*<e��{Y\iq(�&��qS"�3�l�\[5���d�ɽ�*<e�VJUT��� �H4%��&m(���b�{2yiglW�y���9������,(Q'�ƁQu=�U�X��~?�W#m��3+� �?�{�/z��QT�G��J���:ɽ�*<eY[v�_�ɽ�*<eɽ�*<eA��V	{�AJ�EL�cm���fQ�΀�IPd��Qɽ�*<e�Y��2�K+@w�����`�f ��{AQ�OsJɽ�*<eɽ�*<eNM{9q��ɽ�*<eɽ�*<e!�T9�����S����]kKE��ɽ�*<eX��~?�W#m��3+� �?�{�/z�k���C��h
�K=4ɽ�*<eY[v�_�ɽ�*<eɽ�*<e��vVK�`���;�	E\��М}��(H��u�6��/���%��x�#αh�kC�������ʝ�u� <�t-*��h
�K=4����n��rɽ�*<eɽ�*<eɽ�*<e0��葠�Q���Д4��fMT�Ҁ����T�O�4���"#ݷ�x�#αh�kC����J��!㣝˻�%e�܉f��Iă�A����n��rɽ�*<eɽ�*<eɽ�*<eD���p �W"!��ٜ;���D�۳���b\	y`�ɽ�*<e��{Y\iq(�&�� ��E��6��W��#T�.�YС�VJUT���?�(<��ɽ�*<eɽ�*<e��L��	�P�]��cR�o�O�<�ɠ)�Fɽ�*<ex�r%=YF�>���+�5�K��ƐΝ����%�:ɽ�*<e,4���?wɽ�*<eɽ�*<eɽ�*<e7[��İ��u}���ϖ��l�06����b��M&X��~?�W#m��3+� �?�{�/z�k���C�w�	�6�cɽ�*<eY[v�_�ɽ�*<eɽ�*<e��vVK�`^|��]`���G�I�9��p��,ɽ�*<e[��ղ�f� �D�O�h>v����W�����S�ɽ�*<eɽ�*<eҝ[��R�ɽ�*<eɽ�*<eb4�j�[���W��������h���+n�˫Y��2�K+@w�����`�f ��{�>��܎�E#L�@���ɽ�*<eNM{9q��ɽ�*<eɽ�*<e�Gy6+�$�,�IM�+�I頲wD\�w��\��ɽ�*<e�Y��2�K+@w��������
���2�h
�K=4ɽ�*<eɽ�*<eNM{9q��@82�����̟>�ĸ�����d��ve��;�d ���S3b/e�j�!I�2ɽ�*<ex�r%=YF�܎h*�Gm�v[o�I�^ɽ�*<eɽ�*<e,4���?wɽ�*<eɽ�*<eɽ�*<e7[��İ��nꩠ��ʵ&�ӂ[uɽ�*<e����pɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�f#E.��#"�l��Z=�ɽ�*<e�^1�?q�-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\U9��8P�q����d��!I�2�/���%��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc ��9t�������g��h��B,k�׫�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%�)0�/ئ����#m��)/�zC�~��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%���������DC�M���,(Q'�ƁQu=�U�a�磅"��Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���mg��gT�w�W��#T�&ꬶ�Ri=�Z ���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��=�wYh�ǵ��S3b/e�j��T�O�Nd"�O��-&J�� ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡN��Y�T���R���7��$`љR�	���t�nj�'%萚 tɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�f�8��O6@��n�y֜�V��ɾ^1�?q�-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\U9��8P�G��0�@��ɽ�*<e�/���%��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc ��9t����_�av"	;��%���������ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%ז����m�b�!�Z��ɽ�*<e��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%�������~�!8��N��S���ɽ�*<e�+ �0��MK�s�Zɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���mn�W��0^�Lj}��#�˴��56i=�Z ���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��=�wYh�ǵ��nK����Mh}/Y�ɽ�*<e�����l�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡ&H'H�O�%��'X�*��U�������pɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�f#E.��#u���vQ�jɽ�*<e8\(�U�M��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\U9��8P��ܚ���ԯ�f�y��/<��\�T�h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc ��9t������(�-����)P�hx���w�E�@@ZLK|�#ɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%C�k_�pⳮ3f�d]HH��zD��}L�,4��l�ג$OJ�7��D����AP����kP�e�[�[+ɽ�*<eɽ�*<e��x��uۨ�T���]iLɽ�*<e�/���%����qBl�1nmY��
�tx�E�Bxɽ�*<e�/���%����qBl�ڸ�OB���c��LL�cɽ�*<e�/���%�6��j�.QT�'d��!3�_Fɽ�*<e�+ �0�����(T�'d��!3�_Fɽ�*<ea�+Ȳr�s�EŖڿ ˯nkB�J�tx�E�Bxɽ�*<e[a�?~��s�EŖڿ��;�X��d`���N�ɽ�*<e%"	�E׋~\�80R�|�����E_w$[��ڱ�ɽ�*<e7�3]N|���B����(c�lh��-� � x�ɽ�*<e�.���)V���-��Ǔ��x*��@M�aɽ�*<ed��Ję��j<��& �cv�A�ɽ�*<eɽ�*<e�ߐuX�q�&2}��$sN��8H��ɽ�*<e�/���%󬧁��ȉ�id=MK(�b�sN��8H��ɽ�*<e-��)ӕy0�{��NȈ|3k.sb}Hi�X&�M��aO�!�a�+Ȳr���S��$�wyu")�
B�dC�r��ɽ�*<e�U��h��|PZ��9ԁQ�onv>�v��'?�ڷI��bT�>7�3]N|� �#NS)�_Q��'�nL�n삾=Y�Aαh��T�.���)V�ֈ^��}i_Q��'�nL�n삾=Y�Aαh��Td��JęY ]}ړg��ݰI��D��L�𽼛CL��ߐuX�q�N��I-��C= 7\�&~�h����`X#Ԟ����a'�Hs�Ur���2�g�p��bxA��f���ʖ+ �0��0�{��NȈ�e�>��i�p��bxA��f���ʛ�U�ۄ����S��$�w��mf��uВ����E���bT�>�U��h���.z��7�!�қ�Bd:�6�}Zɽ�*<eY�9O=�ʹ�6̴w;��`�:�dnk�/���Z�'[P�u�ɽ�*<eɽ�*<e�
v�ƒm���X��cQ�]�Q�Mɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<eɽ�*<e^��
:�*�~�sh-�ߠwo�	h�[ɽ�*<e[��ղ�f������ܛ�*l�����R��������sk��ҝ[��R�ɽ�*<evS+ё@�˴qZ5�g�}4"{t��HN�E���>Է4X��~?�W#E)�dC��v����W����
���2�h
�K=4ɽ�*<ep<U˸����^1����t��.�-b|X2���H��] �, �W������˾�[(ɽ�*<e1��zfA�kC�����o�2��vc6%8�s���Q�]�Q�M�VJUT���?�(<��ɽ�*<eɽ�*<e�Vz�+#} �h��R�o�O�Nd"�O��ɽ�*<ev���y�1�$W.����|�z ��>��h
�K=4ɽ�*<e,4���?wɽ�*<eɽ�*<eɽ�*<e���,hb��e�d�QWk�HZ�ɽ�*<e1��zfA�kC�����z��=S�w��Rdɽ�*<e�VJUT���?�(<��ɽ�*<eɽ�*<e�]Ӟv��G�I�9��rq��&�c���#�[��ղ�f���;��Y�L����M�L>�;>cc��R��Mbɽ�*<eҝ[��R�ɽ�*<eɽ�*<e��{P���� <�t-*���G�I�9/���?��..+`��[��ղ�f���;��Y�2� ���_d�Ǹ��..
A���ɽ�*<eҝ[��R�ɽ�*<eɽ�*<e���U�&4��%e�܉��+ά���������J�\� R�E��X��~?�W#E)�dC��v����W��Д�٪,EWP���ɽ�*<eY[v�_�ɽ�*<eɽ�*<eA��V	{�A�W��#T���0�7��P�6;7}49�iv (�Y��2�K+׷�����0�堒�c�/���?���h
�K=4ɽ�*<eNM{9q��ɽ�*<eɽ�*<e!�T9�u�P�+H�"hb��e�dB�$Dɽ�*<e1��zfA�kC�����z��=D��M�N�ɽ�*<e�VJUT���?�(<��ɽ�*<eɽ�*<e�]Ӟv�߷G�ey&6��u48ɽ�*<e�/���%�c�i�#J?�{�/z����c��kQ�]�Q�Mɽ�*<e����n��rɽ�*<eɽ�*<eɽ�*<eU�Z�H� �-�!Ɖc�㗟��<�Eɽ�*<ev���y�1�$W.����|�� �"y&�sn5&;�Q�]�Q�M,4���?wɽ�*<eɽ�*<eɽ�*<e�|.���s��@B�#h��4�(T�F(��ɽ�*<ev���y�1�/���>;�#	�q��IX;ɽ�*<eɽ�*<e,4���?wMͿ���q�����&�R@I�K�E���D�M�N�頲wD\�mk��畬�ɽ�*<e�Y��2�K+AC�c�Z�!��pX��ɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<eɽ�*<eșQ�z�~�0/:�,Nv8y�P����g�������$����sbT��82�9��P�6;7}�&ZReX�ɽ�*<eɽ�*<ex�\�uɽ�*<eɽ�*<e+�n�/�G/���?���H�p^|��]`�ɽ�*<e[��ղ�f�oc�v^��J_���Q�]�Q�Mɽ�*<eɽ�*<eҝ[��R�ɽ�*<eɽ�*<em�}�����OG}Db�� �G�\�<��;�sɽ�*<e1��zfAA��y^G��B���b�ɽ�*<eɽ�*<e�VJUT���?�(<��ɽ�*<eɽ�*<e�e��\ȟ)�;C�Q�S3b/e�jɽ�*<eɽ�*<e�����l�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡN��Y�T���/�]� �#hL��>]����pɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�fH����)x��A:!�4�i�9����^1�?q�-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\U9��8Pꔖe�8���!���s�-�/���%��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc ��9t����g�#w�'�S 5l�������ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%Sv(a�iP��%e�܉�j�<�U�q(�B)�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%���������DC�M�jHi��r칌,���+ �0��MK�s�Zɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���m��H�pf�B;i*aކ���jqi=�Z ���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��=�wYh�ǵ�t:�󫓔ɽ�*<eɽ�*<e�����l�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡN��Y�T�z\���ɽ�*<e����pɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e�
O]�S�7�V�B�f܁:ze��d��;}x���ɽ�*<eS�;��$�Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�����/�\U9��8P�S���Γ1��#�s�/���%��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��p�^���Lc ��9t���_tp�n�.]\� R�E�ի�����ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e�MKZ�K������%B}�k���u���vQ�jɽ�*<e��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���/���%���������DC�M��'X�*��U����:�<�.�ؙCB"��,#ɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e���	$���2U���m��G�I�9���(�-����)P�hx�E���G�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��=�wYh�ǵ��YI �_��f�y������&8_K��c��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e[)�i������e6�ڡ����Ve:�X��\��	��F!(�|��\yJ�	;.
�5�ג$OJ�7��D���O�*����J��}�e��e6���Xz2Y2�h^ӽ6���JFV-O�;8W�f��Y��M�]���%����l��^���Q8��;�#��l�,�yU�h^ӽ6��ӸP�[$��fE�ݾa8Z*�h��bo���s�AFqi�3qfVA�0 yɽ�*<e�k�H�� E")��ҜóxW.��ɽ�*<e���m#P�ͮkIR�6������Ue)��fVA�0 y逭R���D�2;LS�?ߐ��&zl��h�ʰC*u�h^ӽ6ԓ����[��WH����/���%�W� �G�+�USm��]²Gװ�u���^!�]q���r�؅��]_��;
鿤ｮ�h4���Yx�.�#d����F����:^���T����ɽ�*<e3��`qP�2��Mc�h4�&�}O��zɽ�*<eO����S�h^ӽ6�O�[d��ɽ�*<e�/���%��r��B #�+�r<5�5H�n�?Y':ɽ�*<e�9��CD�v���Sy1���h�C �G?�L���yFp"Ud����F����:^���b���~��ɽ�*<e+���\�P�R�p�ČO�;8W�fH�T��qKV��G��E")��Ҝo(�;Gx���!�H��(�Eqx�M��I�\�`�P�J��wP��9�ɽ�*<eA�D�/?8�q���n`��r��E�
�*��@M�aɏ@xJ��h^ӽ6�J�k2����J��V2f�/���%��l�{R�F!	�bđxjt�ݯ�ɽ�*<eC�F���ƶ��]_��;�~�c�9hfVA�0 y �n8�]�d����F��� ����~��0�K��ɽ�*<e�Sñ8yY.�n�	10}o<]A�|�ɽ�*<e_�(/�Z�E")��ҜΔ��B��� �G?�L���(�Eqx�'I�5�øxQ@Q�;L	��D2ɽ�*<eӭ0��N����/'�6ɽ�*<eʡB��&yh^ӽ6�bN#D/Qi�W���8���}�i��{c���Ӫ
��
�������%ɽ�*<e{�O����B���Sy1o���R�-�	F��ݏ��������[d����F��#��V�>���u&D`ɽ�*<e��r�����{�h&��v@�.�1 ɽ�*<eB�Q�P�E")��Ҝ�Z��;���ɽ�*<e-��)ӕyd����F�{`is3Z�fVA�0 yɽ�*<ew�����s�.�n�	10�[m5t�ɽ�*<e-&�
:lݲE")��Ҝ��@��[�ɽ�*<e�Fp�AA��j�Tu?4�v9��A�􄘠^!�]qɽ�*<e�ˊ��'�?���n�0ilw|ɽ�*<eT6qRT*nh^ӽ6�����H
�� �G?�L���/���%󬦟�Ly��h���*b���]iLɽ�*<eI?��*�}=�;!���~�L���ɽ�*<e�+ �0��ȩ�h�<L8��=HI~��a�l��ɽ�*<e$Q0��0�{���`�)IjJ�+Rx#5��.�;7�3]N|���}��u�ɽ�*<eɽ�*<e��U�ۄ��	�K�r����nI�CJoX`PV]�/���%�wg�� �� ��C�WaG��ɽ�*<ed��Ję�f�Qu�\ �`Ù�Ÿ�n��
���Wϓ��B�������	H�%1#�,�vL��U�ۄ���!���7�%\�j׸'��^H�/���%�1� ,��"��F�t�e�&�W�Lƍ��OL,4杖�#ڄɽ�*<e1? ��6�+t�c�K�]��s�kɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�-��fΡ��k��4t�pԖ�����Mhɽ�*<e[��ղ�f������ܛ�*l�����R��������sk��ɽ�*<eɽ�*<e�VJUT�����od�t�[.�[��?����w��\��ɽ�*<e�����+���G:fGv���&�;���*������
nP
,����c�´j��B�oO\[5���d��VJUT���?�(<��=K��Hk{��n�v9k��]kKE��ɽ�*<e�Y�3�9��F�t�e�Q��8��y	&-l���P|P�퍓�rlV)iz������$"���y��ɽ�*<eҝ[��R�șQ�z�~�0/:�,Nv8i�e�0ɽ�*<e�Y�3�9��F�t�e�Q��8��y	&-l���P|P�퍓�rlV)iz������$�k|~.�pɽ�*<eҝ[��R�!�T9�G�S$
��!&���S+��������&�JG��b�j��Eh����
lD��#��u��^1�������~���=���Ki���!�)��&ZReX������m�}�����OG}Db�Sv(a�iP�<�ɠ)�Fɽ�*<e�������Br(�&G!1���s�D�<@m̞���&m(��ϑi���8xH��N�ƣw�	�6�cx�\�uɽ�*<eD���p �W����j�D��rq��&�c���#������+���G:fGv���&�;���*������
nP
,����c��c�~Vp�M�L>�;>cS|!kbrB�?�(<���H�خ���v蛍::#E.��#��z�IYLy�q]�iʳ1��@�� ���q|���mVW��c�=��[�sr�G�^6,v��n��g�]C��(ګ���%e�܉�V�� ��ɽ�*<e7[��İ��f�Ӗ�F>���y�a��b\	y`�ɽ�*<e��@�� ���q|���mVW��c�=��[�sr�G�^6,v��n��g���"�[��I<����<{� ̛#ɽ�*<e)_�6-�p�V�*��#��e�8���!���s�-@�j/�j��ڭWH��EZ)eb?S�)��ש0��y�;Xz�����phl���q|����A�c��ԃߔ�B���NM{9q��A��V	{�AJ�EL�cm?����ɕ?kV7�(T�F(�Ś����+���G:fGv���&�;���*������
nP
,����c����'8��Lj}����g���?�(<���t�<=��BDw��?p�H����Q�/ʛ�_�wɽ�*<e��@�� ���q|���mVW��c�=��[�sr�G�^6,v��n��g�J�&M�)j�]��s�k����n��rɽ�*<e	���j�~)�4hK���j�<�U�qɽ�*<e��������:eLE7��\V@���AE
!�ɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uiԙ�&�Vb�m=����9M�(=��49�iv (ɽ�*<e��������:eLE7��\V@��w�	�6�cɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e�#f̨�~��G�=6m�B���ɠ��r\���ֻ'��\yJ�	<�i�~��)G5�td'�b�]���ɽ�*<eɽ�*<eɽ�*<eY[v�_�+�n�/�G�����d<��pR0N���U�'
Rٰ���˫��/���%�\���ֻ'��\yJ�	l\g�Z���<���^��y���C�ɽ�*<eɽ�*<eɽ�*<eY[v�_�+�n�/�G˃�6��Rb��wv�&;���7dɽ�*<e�Y�3�9��F�t�e�&�W�Lƍ3c�3��2@�ࣨSɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�!�T9���	3�Zq��()zӺ_gɽ�*<e�Y�3�9��F�t�e�W���ߺ�i�TF�ۣ��X�Y6�M
����ɽ�*<eɽ�*<eɽ�*<eҝ[��R�X!1e�R�5`��xa�׍hCɽ�*<e�Y�3�9��F�t�e�W���ߺ�i�TF�ۣ}��&�rS�h
�K=4ɽ�*<eɽ�*<eɽ�*<eҝ[��R���������k_�:#_���K�`ɽ�*<e�&�JG��b�j��Ehf�+3yH&�t,�M"�Ž��g�@P,͔�W�7�ɽ�*<eɽ�*<eɽ�*<e�����$Ǟ�2ߊ$�l�	��pw荦xy�cV8��+ Z@�j/�j��ڭWH��3�A�f<㋞�TUn��!`h FH�
�̸B�����y���C�ɽ�*<eɽ�*<eNM{9q��"Rݗ]T��G5�td'�e#<�޼Ũ�^��P#��U��Z@�j/�j��ڭWH��3�A�f<㋞�TUn�ñ�*�jCe�V8��+ Z�h
�K=4ɽ�*<eɽ�*<eNM{9q���m�v�����<���^��Y�Ű�\�kܥ��qɽ�*<e�&�JG��b�j��Ehf�+3yH&�t,�M"�����.�NH�h
�K=4ɽ�*<eɽ�*<eɽ�*<e����옯��U�&4�ҍ�g8��������&ꬶ�R������ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�f�8��O6Nl�>*�2�G���_Db��x���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�����/�\G�P�1�	��=#c?��Z�ØKρ�XcQtp�)�پ������8B`}�FW,P���{Z��
�rt��l�-�b���~��4�1i�Jc2d����F��\	�je�1���b2ޏ� �G?�L��{ �L[�HzdI�4R��z��f��4.�����Sf�H���dd����F��A��~2��fҡ�^��L!�%��+�xՑ*�.�, ������b2ޏ�fVA�0 y�*����*"h^ӽ6��J��}�eC��8�xWf�/���%󬖡���2��
��
����f\�,�ɽ�*<e�u�;�"��]_��;��'g�;S1��<N]��q�����d����F����.ޛXSpL?l�ɽ�*<e�H�i3ﭠO1��	��VZ uD�H�T��q��qz�WE")��Ҝ�P��Ti��a
0�x�(�EqxP��E��ccr�j�����k�:?o
ɽ�*<e{�����Z����bX�ZH�c��ɽ�*<e��P�/�h^ӽ6�%���Nbq,1�Yބ��/���%�6� �����USm��]�fVA�0 yɽ�*<e�(	"<���⥦���G#��Cɽ�*<eT�-5F�nd����F��#��V�C�2w��Z[��!��bKٌ�٦7iJ	���y�j�(��aO�!��d�Տ�E")��Ҝ#"܇a��'~]����(�Eqx�j�Tu?4�\�`�P�J�ܒ��5H�ɽ�*<e[N����br�D�2;L	9��Fgɽ�*<e�
��Y�6�h^ӽ6�>�J#��(ɽ�*<e�/���%�j�Tu?4�:9y����B�p�?�ɽ�*<ex�g� ����bX�Z��A�a�l'ɽ�*<e[a�?~��h^ӽ6�Hk�K{�ԵL	��D2�/���%�j�$�'�Φe�>��9�̖g�%���ɽ�*<e���(�����jx���J���9��ɽ�*<ea�|xd����F�`�� �P1s��^!�]qɽ�*<e�jI�1�;ż��Q��R�k�!�ɽ�*<e��ލk�׫���;��ҟ�d	ɽ�*<es'Syo���<�)3=���K[�k�ɽ�*<eɽ�*<e/q���±�T�y:t�n�5Ǔ��G�tx�E�Bx%"	�E׋u:�`O;�~�T�ȭL���2�-g��H���gXF�+����꣺�X�#e<�P�XB�4M3}���5�l&2}��$sN��8H��ɽ�*<e�.���)VOL$���5�֎%;�#�,�vL�U��h��$�������a?���|\pɽ�*<e-��)ӕy��y����A�O�����'5{��UĖZ�'[P�u�ɽ�*<eɽ�*<eǋ'H)�@w����a���h
�K=4ɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e�4����k���A�X:胮."1Do�ɽ�*<e$����sb����o=�����bC�x���b��6�-4�)�_πZ<�}U�'�:j���+�K�o��c�{��%B{$�"l�+���š�	"�$ɽ�*<e�,��T"��T�����)�堒�c�)u/��L�<Q�]�Q�Mɽ�*<eNM{9q��ɽ�*<e	N�9���� 4���:o�QT�G!���s�-ɽ�*<eO��'��f0%ڡπ�eפm���˾�[(�h
�K=4ɽ�*<e�����ɽ�*<e�Vz�+#} �h��x��[�y��aކ���jqɽ�*<emD�ْ�Ad ݰm�H ��E��6��W��#T�.�YСɽ�*<eҝ[��R�ɽ�*<e��&m�an����g�?�:p׌,㗟��<�Eɽ�*<e�,��T"��T�����)�堒�c�ɕ?kV7�'~_�~Nɽ�*<eNM{9q��ɽ�*<eT��%��G㗟��<�E�4�ҷE��D�j�)Iɽ�*<e�Y��2�K+A�O�����`�f ��{U���g(ɽ�*<eɽ�*<ex�\�uɽ�*<e?������ex���u�P�f>;�݃��������/���%���7�1��kC����J��!㣝��v[o�I�^ɽ�*<e�VJUT���?�(<��ɽ�*<e7[��İ�����э�� ��P�6;7}�~�p[�3�$����sb����o=$W.����|�z ��>���T�O�M
����,4���?wɽ�*<eɽ�*<eD���p �W"!��ٜ;��FZ����Nd"�O��ɽ�*<e�,��T"��T�����)�堒�c�0ڧ�AO4ɽ�*<eɽ�*<eNM{9q��ɽ�*<e���U�&4��C�_@���rq��&�c���#�X��~?�W#��}��N?�{�/z��&�ϔ���2��Aqzɽ�*<e����n��rɽ�*<e+�n�/�G��rq��&�NB�q�vȮ�^q.J1��b��M&�/���%���7�1��kC�����z��=D��M�N�ɽ�*<e�VJUT���?�(<��ɽ�*<e��DO�y4�{fs��.vr(HU�Qɽ�*<e�/���%���7�1��kC�����z��=S�w��Rdɽ�*<e�VJUT���?�(<��ɽ�*<e�٣�eo��T#��Lg��K�am@��wo�	h�[[��ղ�f�2���K,JP�>���"vЅ\��b�]���ɽ�*<eY[v�_�ɽ�*<e�E�$n�d�K�am@�c�ţ�`��Su���eɽ�*<eX��~?�W#��}��N?�{�/z�(��ʸG��h
�K=4ɽ�*<e����n��rɽ�*<e+�n�/�G��`K�f����qNd"�O��ɽ�*<emD�ْ�Ad ݰm�H�LMǊ��..
A���ɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��K��@�BK�K�K�{�!I�2ɽ�*<eX��~?�W#��}��N?�{�/z�:�Y�e��Q�]�Q�Mɽ�*<e����n��rɽ�*<e+�n�/�G�߷G�eyw荦xy�cV8��+ Zɽ�*<eO��'��f0%ڡ�6S�k�=�!�(I���33��0ɽ�*<e�����ɽ�*<e8�q�ѱ�V8��+ Zmm<�=T��d��-QJɽ�*<e	�?�o�.��׈{w�JAv�'�Bɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e�
�Ӛ�.����Ş��i9n��5�ɽ�*<eɽ�*<eD�d�2ud��ٰ#sf��Iă�Aɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�Ef�]�'� ��h/��b��M&ɽ�*<e	�?�o�.��׈{w�J�^ {�Eɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e��Ԫ�N��iAfyl�ދF��ݕٰ���˫��/���%�H'b6]Ȍ���\�m�B���m�����ɽ�*<e�VJUT���?�(<��ɽ�*<eB��gJ��A���4�Qp?0��l�-ǿ�K�am@��wo�	h�[�PI߬H������ȁ�˃�6��Rb��33��0ɽ�*<eɽ�*<eY[v�_�ɽ�*<e��#)ϫ��K�am@�V�D�VO]=,�o��vɽ�*<e�����	Ď����f�[���MĞ��ڭ�oqE�ɽ�*<eɽ�*<e����n��rɽ�*<e+�n�/�G�ƚ�읶���]������ɽ�*<e[��ղ�f�2���K,`E���փ<�~v3����U������h
�K=4Y[v�_�����2(�s:<�\��	3�Zq�B`�M����-��/���%���7�1��kC����m�@�-�F�]��?�`C�..
A����VJUT���?�(<��ɽ�*<e��_NN�ζ���]�؊��SV8��+ Z[��ղ�f�2���K,`E���փ<�~v3�����'����V8��+ Z�iE����nɽ�*<e"`�cd �!�(I�r�++�����/��Z �^���<���^[�Q��S���7�1��kC����m�@�-�F��I�|�ЮH���<���^#z�͌�?�(<��ɽ�*<eD$敃���pR0N6�2��4Y��# N��ɽ�*<emD�ْ�Ad ݰm�Haa24�2G7����^ {�Eɽ�*<eҝ[��R�ɽ�*<e�JLs�����_z+Q4�Q�H�:���:��*ȫY��2�K+A�O�����Sd�~�fT ��w���Av�'�Bɽ�*<ex�\�uG�k`>-:���"��hρ��Ş��i���P�V?��a��{e�ɽ�*<eO��'��f0%ڡШ6�E���hƁ�,f��Iă�Aɽ�*<e�����ɽ�*<e�Ef�]��_z+Q4�QPn���&���!�(I켥����TUA�O�����Sd�~�fT ��w���"�#F��8����T�x�\�uɽ�*<e"Rݗ]T��G5�td'�e#<�޼ń��P�V?8����		%�����ofO��'��f0%ڡШ6�E���f�M�
V8��+ Z�h
�K=4�����ɽ�*<e�e	�5S�B���@%He�����E�����ɽ�*<e�,��T"��T�����)yyֶ�T@E%��D�&�y�����ɽ�*<eNM{9q��ɽ�*<e���P��r"L�ń|%<R|=-�z�`u�tu1�D@u{�l�ʶ���u�[��$�ss]d��9�^8�7ɽ�*<e����n��rp�^(]e���}��h����`K�f8l��	�%Y�g�E�����P�dE�0(|�:B�2ƍ�zC�'��������v믜�LQ�]�Q�Mɽ�*<eҝ[��R�ɽ�*<e��K��@���>�dS@<R|=-�n �u�HYaU�.n��p�l�ʶ���u�[��8�����}�\U�>:�ɽ�*<e����n��rɽ�*<e+�n�/�G�߷G�eyp�^(]e����j�M�}�-��%��ɏu��7)��S�c�Y�=��<�wj@�ɽ�*<eɽ�*<e�����ɽ�*<e�����i���}hc�f���9TI���.�NH�Y��2�K+A�O�����Sd�~�fT�[V�`��,\�8� 'z��9�^8�7x�\�up�^(]e��#ӛvn�J���Ş��ip�^(]e��#J�����`����-�O��'��f0%ڡ��㟰��TM�B"�OVQPXp�P�Q�]�Q�M�����ɽ�*<e�Ef�]����}hc�f���9TI�����7�Y��2�K+A�O�����Sd�~�fT�[V�`���S�)n%�\U�>:�x�\�uɽ�*<e��Ԫ�N��{fs��.v2X0u0�pM*��U����/���%���U�?��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT��ȅ5�+�!m>��e6�ڡ�h�&u��p)2���@�h2uvÐ�2@�3�#[���HK
ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��p�^���Lc �v�l������4\���鳣���`��V�,�W]�ͻlU�� <�ZBg�cG4�NP�g���=z Ҡ�z;���ӷ�l2.��k���-F��lB��dzMp/�ar��\R`S�5�{AM�ɽ�*<e���[��c��#�����	/���U�ۄ���d���/)��H/��ɽ�*<ed��Ję���'�D&����A��tO�4�!���7�%�&�����V����Fd��Jęf5-�M0,�3��x�K���tO�4�!���7�%$�A��˼���d��Ję4��Wzhp�I�ۿww�佦i0Oh�!���7�%1�@ͫ�����e�ʝd��Jęs�Ϭ(�����Z){Q��r��<�-<���� �2���K,`E���փ<�t�jA(OZ�'[P�u�ɽ�*<ew�;L�::=�Y��r����&6ɽ�*<eɽ�*<eɽ�*<e,4���?w:j���+�oaf�	��,��/�=X]ɽ�*<e�Y��2�K+��Qݓ˟s4�)�_π ����������'�e����ǄA�8���K�o��c�{��%B{$���}���49�iv (�Y��2�K+A�O�����Sd�~�fT ��w���^ {�Eɽ�*<ex�\�u�&�|�D�#f̨�~a��#;�Nd"�O��[��ղ�f�2���K,ݥ D���z}x���Q��AE
!�ɽ�*<eY[v�_�+�n�/�G���q��l2`�
��(yaf��ٿ[��ղ�f�2���K,ݥ D���z}x���Q�W:�=����ɽ�*<eY[v�_�+�n�/�G��`K�f࣏�>�m�B���D���&�K2���K,ݥ D���z}x���Q������d<��5�2-Y[v�_�+�n�/�G�����d<��pR0N���M���ٰ���˫�[��ղ�f�2���K,ݥ D���z}x���Q�˃�6��Rb��33��0Y[v�_�+�n�/�G˃�6��Rb�y��k~�f��S�Hɽ�*<emD�ْ�Ad ݰm�Haa24�2G7����^ {�Eɽ�*<eҝ[��R�\/l�<�]��<}�l=2���mɽ�*<eO��'��f0%ڡZm��B��H�@�p1�AE
!�ɽ�*<e�����H�*��h�Aa���d1�W�D6�fɽ�*<eO��'��f0%ڡZm��B��H�@�p1W:�=����ɽ�*<e����옯��U�&4�h^�!�����ym��Aٰ���˫�O��'��f0%ڡZm��B��H�@�p1�����d<��5�2-�����w[i����Ç̸B�����\>�_�V��P �޸����ofO��'��f0%ڡZm��B��H�@�p1˃�6��Rb��33��0���������Ħ�
V8��+ Z)�[��w��\���:�<�.�ؙCB"��,#ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곑f�[��!Nd"�O����{��Q�h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ��`���)6�-�@v�ɽ�*<e-&J�� ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�f�б�͞8;7v��������pɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�����/�\U9��8P�6���N%��|�/��=1��[>�V�/eJR�k�/eJR�k�/eJR�k�,q'�Q�OQ�]�Q�M��M�R��Lc �Ij�a�*c�&�c���	����K��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���	D��:�^�����%��j��\�P�}7"\]e����,Wɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<ej	�%w\�����R��kq6v��%`���ɽ�*<e(�B)�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eu;�Qݷ�2U���m��̲�E6�y�k">z��a�磅"��Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곛�y�v|�iP��[P��{��Q�h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ��|�KLǍ�V����2ɽ�*<e�����l�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�f''�����J�J=���	���t�nj�'%萚 tɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�����/�\U9��8P�)�7h����X���W�
U�K;ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��M�R��Lc �v�l��Vh��S�zC��YB�gN2E[5���ԉ[��Q�)yӡ'�7�e�SuJg��/.�w <>k��h4�����#}w|�)�S�^5d�<l]j^a5k:e�."�v���l^��V���@}tV��^���>�A*��O2�9�L>2�kΟ���T�u�5�808;lAf ��)��v���l^�M��I�cr�j���[���K��ɽ�*<e)G;�?��I.�, ������b2ޏ� �G?�L����:Tǃ�h^ӽ6��IuW�������/���%�DY��x�v���f�9�O�����ɽ�*<e�jQK�6�	�y���:�S�Z�:���B�p�?� }�U�Pyd����F����.ޛ���1��ɽ�*<e�V/�P�R�p�Č�4�d���ɽ�*<e�Ewp��IE")��Ҝ�P��Ti��<��y�(�EqxP��E��c�"�YZR 6�q��ɽ�*<e��S�NW�ʵ��bX�ZE^�X,6�ɽ�*<e�Д��ʝh^ӽ6�Έ��"�q�ɽ�*<e�/���%��Y�Dxu��USm��]� �G?�L��ɽ�*<e1���\#����Sy1"�#$W&��L�0S0�?��<d����F��#��V�>Ey�U#�ɽ�*<e��$P/R�7iJ	��C�^a��ɽ�*<eyu��}��E")��Ҝu���|�����~M�D�(�Eqx�5D@/V��6�����L	��D2ɽ�*<e�;"���3r�D�2;LF�
('f�ɽ�*<e�U��h��E")��Ҝ � 	��#�ɽ�*<eL�@t�Z�s��V���@}:9y���}Mw�Ψɽ�*<e^iB�j�f��O�D d�4Oq��ɽ�*<e�k��)�h^ӽ6�Hk�K{�ԵH�T��q�/���%�S��\a�Z��p�q�xU�ީ�Lɽ�*<e� �;�m���jx���JMWK5�ޭ ɽ�*<ef�R�X6�Vd����F���'?�ڷI�tx�E�Bxɽ�*<e1M ҵ��[��^Us&�'2g�Doɽ�*<e%{5��0 ���Kx�?�^*���ɽ�*<e�v���l^N���Ir�nO9���c��LL�cɽ�*<e$Q0��0�{���`�)IjJ�+Rx��>�G�@7�3]N|��|���A��_�4��(���`�2]��tO�4�!���7�%fKˍʔ��	kU�f�Z�/���%󬧁��ȉ�id=MK(�b�sN��8H��ɽ�*<ed��Ję�� �2�ہ�-���ɽ�*<eY�9O=�.XҎ�~Sx=��/K��#�����Xv�kɽ�*<eɽ�*<eg��1-P��V]��%�ɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<��G�x9��FE�&I��}Kg��@հɽ�*<eɽ�*<emD�ْ�dh89QN��hz�;3��PY���F��
�W���[�&`�ժH��������L���xr��<I}����hd�m��"�,w#ɽ�*<e�Y��2�K+ҫ�0�7�v����W����
���2�h
�K=4ɽ�*<eY[v�_�ɽ�*<e5�?��
��;�d ��Hk�P��|�W����sp�ɽ�*<e��w�&��^Sx=��/π�eפm���˾�[(�h
�K=4ɽ�*<e�����ɽ�*<e�Vz�+#} �h��x��[�y��aކ���jqɽ�*<e��w�&��^Sx=��/5�d��X,��b\	y`��h
�K=4ɽ�*<e�����ɽ�*<e��L��	�P�]��c�����U�:���y��Vɽ�*<e��w�&��^Sx=��/�ч�t}�,�IM�+�IQOB-�y�ɽ�*<e�����ɽ�*<e���|���(zSȢ�|N)�/Ԁ;�DhY��F�ɽ�*<e�l�FD�V��jU�.x���Y.w���`2���ɽ�*<eɽ�*<eҝ[��R�ɽ�*<eIh�����jKfz=�8;7v����ɽ�*<e�Y��2�K+ҫ�0�7�v����W���P�6;7}�&ZReX�ɽ�*<eY[v�_�ɽ�*<e!�T9�u�P�+H�"��FZ���ͻ�%e�܉�j�<�U�q�l�FD�V��jU�.2� ���_d�Ǹ��..
A���ɽ�*<eҝ[��R�ɽ�*<e��]/߷�W��T�O��C�_@�"�d�;�ɽ�*<eX��~?�W#-KB�i�`�f ��{AQ�OsJɽ�*<eɽ�*<ex�\�uɽ�*<e�H��g�2$��Z�!�I����!�r칌,���/���%󬷌�{�}f$W.����|�.k-���!Eg2�����Q�]�Q�M,4���?wɽ�*<eɽ�*<e0��葠�Q���Д4��k���C��!I�2ɽ�*<e����^��kC�����z��=D��M�N�ɽ�*<e�VJUT���?�(<��ɽ�*<e��DO�y4�{fs��.vr(HU�Qɽ�*<e�/���%󬷌�{�}f$W.����|̃��h�&,.�YСɽ�*<e,4���?wɽ�*<eɽ�*<e�����I��rH�&V8��+ Zɽ�*<e�l�FD�V��jU�.+[�&�����<���^��y���C�ɽ�*<eҝ[��R�ɽ�*<e��{��s����4�Qp?�*���U ��:��*�ɽ�*<e[��ղ�f�!��QE����~��!W:�=����ɽ�*<eɽ�*<eNM{9q��ɽ�*<e���U�&4�h��4��lR����P�ɽ�*<e$����sb�F{N.J?�{�/z�v�7�w��h
�K=4ɽ�*<e����n��rɽ�*<e+�n�/�G���q���&�M���ɽ�*<eɽ�*<e��w�&��^Sx=��/�:�W�Ӡ��\U�>:�ɽ�*<eɽ�*<e�����ɽ�*<e�� Qx����H�3���!�(I켔-�э�g�[��ղ�f�!��QE����~��!�����d<��5�2-ɽ�*<eNM{9q��ɽ�*<ew[i����Ç̸B���7)�ĝfһ\�kܥ��qɽ�*<ew�;L�::{���	�����c�h+�0�ɽ�*<eɽ�*<e����n��rɽ�*<e�N*z+N����`K�f�"���Nd"�O��ɽ�*<e=�i>�N���0yB�̴VQPXp�P�Q�]�Q�Mɽ�*<eɽ�*<e�����ɽ�*<e�Ef�]�'� ��h/��b��M&ɽ�*<e	�?�o�.�	c�W.�ҽ�0���Ѓ��&ZReX�ɽ�*<eɽ�*<eY[v�_�ɽ�*<e���������f�fQI �"�#F��8#��U��Zw�;L�::{���	��?� :�f|G5�td'�b�]���ɽ�*<e����n��rɽ�*<e+�n�/�G�����d<��pR0N���U�'
Rٰ���˫�ɽ�*<e=�i>�N���0yB�̴���v��{�5�2-ɽ�*<eɽ�*<e�����ɽ�*<e�e	�5S�B���@%fzA?���B�"���ɽ�*<e�F`��� ^ .=2�����g�@P,͔�W�7�ɽ�*<eɽ�*<eҝ[��R�ɽ�*<e
�'63��ׇ�f���@
���B��d��-QJ�/���%󬷌�{�}f$W.����|�o�K��o�G�e�2� ���9�^8�7,4���?wɽ�*<e��*�M��嫑�$�*�q\+m"���~`��rɽ�*<e�l�FD�V��jU�.aa24�2G7����ᦲc�ɽ�*<eҝ[��R�ɽ�*<e��K��@��\�L{���c�XO�_ag�̸B���%��Й�-KB�i�Sd�~�fT^�0��ş{M�y0��bm�B���*c�n��&ɽ�*<e"Rݗ]T��G5�td'�e#<�޼ů5�MP��˃�6��Rb�-�э�g�����^��kC����m�@�-�F��I�|�ЮH���<���^#z�͌�?�(<��ɽ�*<eD$敃���pR0N6�2��4Y��# N��ɽ�*<e��w�&��^Sx=��/Zm��B��H�@�p1w�	�6�cɽ�*<e�����ɽ�*<e�� Qx���}&��׶�}.8��lj&��1��[��ղ�f�!��QE��yyֶ�T@ÙEǛ'�h+�0�ɽ�*<eNM{9q���5��[1gԟ��R����HB����}x���Q�..+`��$����sb�F{N.J?�{�/z����P�V?禺��zQ�]�Q�M����n��rɽ�*<e+�n�/�G���q��nL����a3��|��V8��+ Z��w�&��^Sx=��/Ш6�E��R�a�G��̸B�����y���C������ɽ�*<e8�q�ѱ�V8��+ Z�_z+Q4�Q~��/��K�am@�dZ��`R�$ҫ�0�7�ݥ D���z}x���Q�˃�6��Rb��33��0Y[v�_�ɽ�*<e��#)ϫ��K�am@����}2�K�E%��D�&��b��M&X��~?�W#-KB�i�Sd�~�fT ��w���^ {�Eɽ�*<ex�\�uɽ�*<e��Ԫ�N�Ml��+aC~�[V�`��G	�ģ�BH���N��g�����6��o����a��ר�d��2��.ău�Y�',4���?w����M�%Y�g�E����$�*?Ѳչ���7Ց�X2��~`��r\_*X�#~v'�w�֬����K��NJ��� ..
A���ɽ�*<eҝ[��R�ɽ�*<e��K��@���>�dS@<R|=-�n �u�HYaU�.n��p�l�ʶ���u�[����Ķ���U2�1D���ɽ�*<ex�\�uɽ�*<e��Ԫ�N�Ml��+aC~�[V�`�����@��=�$�⥴F�1g�����6��o����a��רO4����U�b9v�B	�,4���?wɽ�*<eɽ�*<eM�Uy-V9?Ѳչ��&�����ڧ\�kܥ��q�l�FD�V��jU�./��+�ͼ�f���9TI���.�NH�h
�K=4��۩�f6<<R|=-��]2�f r�S�D�<R|=-��X�Y6������5C-KB�i�Sd�~�fT�[V�`��zǙ�7��h��x�\�uɽ�*<eW���P�#��6*+�'p�^(]e��A ��%��b��M&����^��kC����^��N2�{�&�����ڧ�^ {�E�VJUT���?�(<��ɽ�*<e:��8*$7��WG��Kгj����N0ɽ�*<e8\(�U�M��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�����/�\U9��8P�k���C�\#����r�..+`��K��c��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT��ȅ5�+�!m>��e6�ڡ����Ve:�X��\��g�����6��n��_Lq f�&�������Y���:cl ��C��z󚅔��Q}���5�lcnNMG���뿓�؋��Ŵ�����e��Ċ�|�J���ɽ�*<e��pJ�1�7�A�7e���5�-��)ӕyƛ�R�n�8s6��ZL	��D2�.���)V��w�o傏(�Q3X,�+ �0��L��P�a��M�G�1�2Zs��Q,��.���)V�GT��)��S����{�+ �0��L��P�a��t�W����_����mQ��.���)V�yA�ߠ��j�;�y	�L�q�_�L��P�a�ĭ��l���v�����R���.���)V��|�������	z�i�j��lp���O��y����ҫ�0�7�`E���փ<�t�jA(OZ�'[P�u�ɽ�*<ew�;L�::=�Y��r����&6ɽ�*<eɽ�*<eɽ�*<e����n��r�G�x9��FE�&I��}Kg��@հɽ�*<e[��ղ�f������ܛ�*l�����R��������sk��ӈ����
%:�=~<���%�6��Aiq��%ɽ�*<e�l�FD�V��jU�.Z�?�v&i5%�u�){K�\U�>:�ɽ�*<eҝ[��R�!��2����jN�̓������P�ɽ�*<e����^��kC����K��H7Mc(J ��M
�����VJUT���?�(<���K��@�G5��3iv�Su���e�/���%󬷌�{�}f$W.����|�TErǃ+�\�r+�=��h
�K=4,4���?wɽ�*<e��t5��;LӚٿr-�G5�td'� =��jB��F{N.J?�{�/z����P�V?� �^J��yϦM�|.{� ̛#ɽ�*<eB��gJ��A���4�Qp?��&�E@s��K�am@��m9C?'n�-KB�i�Sd�~�fT ��w����"vЅ\��b�]���x�\�uɽ�*<eن�\�)�e#<�޼ż�l�G��ɽ�*<e�l�FD�V��jU�.aa24�2G7����^ {�Eɽ�*<eҝ[��R�\/l�<�]��<}�l=2���mɽ�*<e����^��kC����m�@�-�F�]��?�`C�..
A����VJUT���?�(<���K��@��@��\�kܥ��q�/���%󬷌�{�}f$W.����|�o�K��o�G�e�2� ���9�^8�7,4���?wɽ�*<e��t5��;��̲�E6������d<��#������F{N.J?�{�/z���"o��D j��c�̸B���^0�\<efɽ�*<eB��gJ��A���4�Qp?��^� |����<���^�%��Й�-KB�i�Sd�~�fT^�0��ştseQ,�yϦM�|.9�<7���ɽ�*<eن�\�)�e#<�޼ŝ� �v��(T�F(��8\(�U�M��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<eu;�Qݷ�2U���m)�[��"�d�;��+ �0��MK�s�Zɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�����/�\U9��8P�6���N%�&ꬶ�RS�;��$�Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<eu;�Qݷ�2U���m)�[��/���?��a�磅"��Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�����/�\U9��8P�6���N%��|�/��=1��[>�V�/eJR�k�/eJR�k�/eJR�k�,q'�Q�OQ�]�Q�Mu;�Qݷ�2U���m�?ŸAl�6Zg��7��~�,�~Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�����/�\U9��8P�|�� ����!i�#%}ʔʵ�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eu;�Qݷ�2U���m��Moi��vΦ�-C��z�+ �0��MK�s�Zɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�����/�\U9��8P�ɉj�]�!�(yaf��ٿ�^1�?q�-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eu;�Qݷ�2U���m��Moi��v��МB\'��+ �0��MK�s�Zɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�����/�\U9��8P��/1lG%iP��[P�^1�?q�-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eu;�Qݷ�2U���m�|6*]�&��Jd�q/ݖ+ �0��MK�s�Zɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�����/�\U9��8P�)�7h����X���W�
U�K;ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eu;�Qݷ�2U���m�  ƿzp��'a�y�鍕D�3�/j�u�x��b��i���sX!�摠Z����\	�je�1���b2ޏ�fVA�0 yH�5��P�{Z��
�rt��l�-Z���Kza ׺{G��2d����F��A��~2��fҡ�^���%w��v�ߣ��}إ"zdI�4R��z��f��4.� *=5[0�Y�j�9Dd����F����:^���b���~��ɽ�*<e+���\�P�R�p�ČO�;8W�fH�T��qKV��G��E")��Ҝ����2�1��Eݤ/�(�Eqxk�քM5�j�:K�i��t���J}E�ɽ�*<e�l�Y�m��"�  v�C �7�fVA�0 y��xO&��h^ӽ6�J�k2����lg�f'%�/���%������H�ި}E](��^�����ɽ�*<eC�`�� ��]_��;�~�c�9h �G?�L�� �n8�]�d����F����:94�Pz��2��ɽ�*<e%���b`
_.�n�	10]�pTWɽ�*<e�:|�l��eE")��Ҝ�=�_�OU�ɽ�*<eu7���NP��E��cøxQ@Q�;H�T��qɽ�*<e������2�9�F�c����������撗wA�f��h^ӽ6�`q��Z�@T�R��n�/���%�@!!���
��
���-S��N�	ɽ�*<e����:�ـ��Sy1��T'ig���aO�!�M$�mVed����F�}D�4iɽ�*<eɽ�*<e��R�/�x{�h&��vP�5wu��ɽ�*<e7�3]N|���]_��;��Ox�nQ&ɽ�*<e.��x�y�Nd����F�{`is3Z� �G?�L��ɽ�*<e�A����חl-�^�� �xU�ީ�Lɽ�*<e�1q6�\
E")��ҜY;������ɽ�*<e���m#P��P��E��c� Nb '�B��K�ɽ�*<e���Pz%w�?���n���@� �ɽ�*<e��mp�n�h^ӽ6ԥ~3?7`����]iL�/���%�pP3�am���hAU6]?���,	4ɽ�*<e�#wƇv���C�g�{��tr��ɽ�*<e/�WA�Y0�{��NȈ�^�hq>Q��a�l��ɽ�*<e�%������En�]H��Q1���LHH0��.���)V�0�z���m��h{��6.b���ݵYi��Lw�羈�g���.�Dz�.�-��)ӕyL��P�a��$���$t�_rw���+ɽ�*<e�ߐuX�q�oL�P{�Pw\!h��m\ɽ�*<erP/�ۻ�dFK��Z
�i(�?K��#�����Xv�kɽ�*<eɽ�*<eg��1-P��V]��%�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����:j���+�oaf�	��,��/�=X]ɽ�*<eɽ�*<e�,��T"���`χ�a$����^�M�"�ds��R��6G�2���-l	*vNM{9q����;��R�˴qZ5�����9u���
���2ɽ�*<e$����sb�����x�$W.����|txG�z��h'~_�~Nɽ�*<e,4���?wɽ�*<e�Ja�f�ل�%�>v;�jT��_��J�EL�cm�wo�	h�[�Y��2�K+)�ߙmit�`�f ��{�A�c��ԃߔ�B���ɽ�*<ex�\�uɽ�*<eA��V	{�AJ�EL�cm��;�����g�#w�'�S 5l�X��~?�W#
j���?�{�/z�wM�.�����$�c>y�Dɽ�*<e����n��rɽ�*<e+�n�/�G���g�#ww@&T.�f������h���+n��$����sb�����x�$W.����|�� �"y&�sn5&;�Q�]�Q�M,4���?wɽ�*<eɽ�*<e���#B? ��T�i��6s��}�ɽ�*<eɽ�*<eO��'Z
�i(�?��8�z4ؓ���+4�ɽ�*<eɽ�*<e�����ɽ�*<e�h�z��qc�w�LV�/�5�'��,��ɽ�*<e[��ղ�f�}%^Y[�\Vv����W���P�6;7}�&ZReX�ɽ�*<eY[v�_�ɽ�*<e!�T9�u�P�+H�"��FZ���ͻ�%e�܉�j�<�U�q�,��T"�˺-H嵰. �堒�c�/���?���AE
!�ɽ�*<eNM{9q��ɽ�*<e���U�&4��%e�܉�0����P��IPd��Qɽ�*<e$����sb�����x�$W.����|�z ��>��h
�K=4ɽ�*<e,4���?wɽ�*<eɽ�*<eM��u�^8:㋞f����(H��u�6�ɽ�*<emD�ْ�A�^_p�xL����M�L>�;>cc��R��Mbɽ�*<eҝ[��R�ɽ�*<e�H�خ���v蛍::���x4��B�$Dɽ�*<e[��ղ�f�}%^Y[�\Vv����W�!&���S+�\U�>:�ɽ�*<eY[v�_�ɽ�*<eșQ�z�~���;=6
����x4���QWk�HZ�ɽ�*<e[��ղ�f�}%^Y[�\Vv����W�"���y��ɽ�*<eɽ�*<eY[v�_�ɽ�*<eșQ�z�~�к���@��9��I������of�/���%�Iή�%`��kC�����<-`__�V8��+ Z�h
�K=4�VJUT���?�(<��vS+ё@�v�D�,��pR0N����Y�(yaf��ٿɽ�*<emD�ْ�A�^_p�x�#ڴ-P�h+�0�ɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��]/߷�W����G"l..+`��ɽ�*<eX��~?�W#
j���?�{�/z�v�7�w��h
�K=4ɽ�*<e����n��rɽ�*<e+�n�/�G���q���&�M���ɽ�*<eɽ�*<emD�ْ�A�^_p�x�,�)7�1��y�����ɽ�*<eɽ�*<eҝ[��R�ɽ�*<e�JLs����
�Y�7f�OG5�td'�a�k|jZ��Y��2�K+)�ߙmit��Sd�~�fTދF��ݕyϦM�|.Q�]�Q�Mx�\�uɽ�*<e"Rݗ]T��G5�td'�e#<�޼�s$w�h�'ɽ�*<eɽ�*<eD�d�2uc�A�`P�Av�'�Bɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e��eZ�L�G��b�`�Ҧ���-�ɽ�*<e	�?�o�.����n�d��ٰ#sf��Iă�Aɽ�*<eɽ�*<ex�\�uɽ�*<eW���P�#��6*+�'n�E-��bɽ�*<eɽ�*<eD�d�2uc�A�`Pꞡ^ {�Eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�� Qx��ӂ�c�H���!�(I켔-�э�g؀PI߬H���S�B���kȌ���\�m�B���m�����ɽ�*<eY[v�_�ɽ�*<e"`�cd �!�(I���wv�&��9��I������of�/���%�H'b6]�@c}�b�˃�6��Rb��33��0ɽ�*<e�VJUT���?�(<��ɽ�*<eD$敃���pR0N���ᇴM��X���ɽ�*<e=�i>�N� PزK`Q[���MĞ��ڭ�oqE�ɽ�*<eɽ�*<eҝ[��R�ɽ�*<e
�'63��ׇ�f���@
���B��d��-QJ�/���%�Iή�%`��kC����m�@�-�F��9�:~���h+�0��VJUT���?�(<��^�u������h��j�����]� b��ɽ�*<e[��ղ�f�}%^Y[�\V`E���փ<�~v3��>|
ϒ����h
�K=4Y[v�_�ɽ�*<e�`���{R�5`�����P2��G5�td'J3�W�`>+Iή�%`��kC����m�@�-�F�4�)�*�z�G5�td'��C�	�?�(<��ɽ�*<eB��gJ��A���4�Qp?����]6vZ�%�M#��U��Z[��ղ�f�}%^Y[�\V`E���փ<�~v3��G������r����T�Y[v�_�ɽ�*<e��#)ϫ��K�am@����}2�K�n �u�HY49�iv (X��~?�W#
j���?�{�/z���"o��D�2nq�Ř��&ZReX�����n��rɽ�*<e+�n�/�G�߷G�ey���P�V?TO�Ɩ�tzɽ�*<eO��'Z
�i(�?Ш6�E�.8��l@�ࣨSɽ�*<e������B֊ ��f�̚νEn�_z+Q4�Q�m�3'k:��q]�iʳ1�Y��2�K+)�ߙmit��Sd�~�fT ��w����ᦲc�ɽ�*<ex�\�uɽ�*<eW���P�#��6*+�'���P�V?� �^J��ٰ���˫�O��'Z
�i(�?Ш6�E��R�a�G��̸B�����y���C������ɽ�*<e8�q�ѱ�V8��+ Z�_z+Q4�Q~��/��K�am@�dZ��`R�$)�ߙmit��Sd�~�fT ��w����"vЅ\��b�]���x�\�uɽ�*<e�m�v�����<���^�d=�#�<d}x���Q��!I�2$����sb�����x�$W.����|�TErǃ+W=CՂ�z�Q�]�Q�M,4���?wɽ�*<eɽ�*<e�#f̨�~8l��	�%Y�g�E�\�kܥ��qdE�0(|�:B�2ƍ�zC�����y*$�ss]d��9�^8�7ɽ�*<e�	��l\�f���9TI2�h	�r�S�D�<R|=-}!�Lڜh�8FP�G�l�ʶ���u�[��� �ڄ��v믜�LQ�]�Q�M����n��rɽ�*<e+�n�/�G���q��8l��	�%Y�g�E�Y��# N��dE�0(|�:B�2ƍ�zC�����y*8�����}�\U�>:�ɽ�*<eҝ[��R�ɽ�*<e�JLs�������}hc�f���9TI�&!�r8�E�7��Ala�v2}&�PZ�n.{{LZ�"""���<�wj@�ɽ�*<ex�\�uɽ�*<e�m�v����>Ѷe%Ap�^(]e��C�]�Nf�ݏd��-QJO��'Z
�i(�?��㟰��TM�B"�OxL5�M�k/Q�]�Q�M��fT�u|f���9TI�9�k��˅��}hc�f���9TI��~-y7�Y��2�K+)�ߙmit��Sd�~�fT�[V�`��zǙ�7��h��x�\�uɽ�*<eW���P�#��6*+�'p�^(]e��A ��%��b��M&O��'Z
�i(�?��㟰��TM�B"�O2�ia�s�aɽ�*<e�����ɽ�*<e�� Qx��ӵw�LV�/�u���vQ�jɽ�*<e�>1�"@�q26�\�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_��MKZ�K������%��S�b��L{���V݅Ϗm�/
S�;��$�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q����=�wY�@o��W������&�5�D���z���'呝]A���C��&���Q�)y����-���F�ud�^jN�z/32�
���Wϓ���cp��RJlJ���ܡVx��a�l�/��/�8�0qe��]��c=���DХ�Oq�c�]�h�,�B��)��\|}�d��Ję���.���L��+�
��U�ۄ���!���7�%� Q��5ɽ�*<e�%�G��o�d�BjZ@L�cs���U�ۄ�����K�u�	H /�)w$[��ڱ��%�G����A�I�򄷘x������C�I��!���7�%0_S�do5���d��Jęs�Ϭ(�����C�K�e��	�!���7�%1�@ͫ����5)"�0��8����Iή�%`��kC����m�@�-�F�&�U �H����Xv�kɽ�*<e��+�J^�Q��	�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q���4����k���A�X:胮."1Do�ɽ�*<eO��'��P�n�/ͻ�:||hy�6"pUw�����I�� �pQ��/�%×�˴qZ5���,�Y��# N��ɽ�*<eO��'Z
�i(�?Ш6�E�SD+�?M��&ZReX�ɽ�*<e�����㵫�*�	�Z|[s%�o..+`���/���%�Iή�%`��kC����K��H7Mc(J ��M
�����VJUT���?�(<���K��@�G5��3iv�Su���e�/���%�Iή�%`��kC����K��H7�g'P��Său�Y�'�VJUT���?�(<����]/߷�W�LG�������d<�- �Ƈ���Iή�%`��kC����K��H7Z�j"�nm�B���(�ZZZ���?�(<��g*D����Vm�B�����V���/�˃�6��Rb9k/�i���Iή�%`��kC����K��H7�B5+o=�yϦM�|.��ZXd�"?�(<��P�ay��b���4�Qp?wb۳.��:��b��M&X��~?�W#
j���?�{�/z���"o��D�2nq�Ř��&ZReX�����n��r���&B��G��θ��x�H�q]�iʳ1�Y��2�K+)�ߙmit��Sd�~�fT^�0��ş91��?��M
����x�\�uɽ�*<e�m=����9í�>0\͟�:��*ȫY��2�K+)�ߙmit��Sd�~�fT^�0��şAwo��o�ău�Y�'x�\�uɽ�*<e���$�*��́��>��!�(I켥����TU)�ߙmit��Sd�~�fT^�0��ş{M�y0��bm�B���*c�n��&ɽ�*<e����o���S�B���@%;�� ����K�am@�dZ��`R�$)�ߙmit��Sd�~�fT^�0��ştseQ,�yϦM�|.9�<7���ɽ�*<eن�\�)�e#<�޼ŝ� �v��(T�F(��8\(�U�M��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��M�R��Lc ��M��C�IPd��Q�/���%�ȣleg�׿ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���	D��:�^�����%e�2���QWk�HZܓ��z:�-q26�\�ɽ�*<eɽ�*<eɽ�*<eɽ�*<ej	�%w\������~�W%8n�Y��]��J��b��M&��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eu;�Qݷ�2U���m)�[��i���!�)�!���rv�J3�tM/eJR�k�/eJR�k�/eJR�k�_�p�fh+�,4���?w��=�wYh�ǵ�n���k��d.e�&�ͮ�7��fc�Pɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡJR�^��hX�Wk�k�s����Od�����l�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�f?�
��#&'ZC��	���t�nj�'%萚 tɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�����/�\U9��8P�ɉj�]�!�(yaf��ٿ�^1�?q�-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��M�R��Lc �<gcp2��}�-��%��/���%�ȣleg�׿ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���	D��:�^�����%����AYe�u�d}l������ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<ej	�%w\�����R��kq6vc���ġ[��%�w/(�B)�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eu;�Qݷ�2U���m��̲�E6�,�o��va�磅"��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wY�@o��W������&�5G���0��Jf�x�\("��	�wR"]�ͻlU�� <�ZBg)�S�^5d�<l]j^a[���K���v���l^P��E��cSuJg��/.�w <>k��h����8��G�T�u�5�808;l>��J$�~�v���l^�'I�5�tV��^���>�A*�Ӭ��g0��@�D�b��]_��;.�w <>k��h4���5<�����d����F����:^��Z���Kzaɽ�*<e�?is���ئ7iJ	��qz�v�;ɽ�*<e=���5|+E")��Ҝ�}�9��F�Q�)(�Vx���m#P�͓�V���@}���tgv
�!#�Bw�ɽ�*<e�h����"�  v�C �7� �G?�L��zG��.�h^ӽ6ԓ܌���/%X@�S%�/���%�����t\�M�ި}E](�N��ɽ�*<eC�`�� ��]_��;�E�I6�L	��D2d��8���d����F����:94gإ���٣ɽ�*<e���a��N߬�:ǄA�hǳ�o�ɽ�*<e�]��Q��E")��Ҝ:���RTɽ�*<eL�@t�Z�s�kIR�\�`�P�J��b~*R�R�zr��A�lԃ��G�w9�F�c@�8�!5�/�w�Yݿ��h^ӽ6Զ�����֋R��D���/���%��.����G�
��
�����$S�ƾɽ�*<e�\�]�#����jx���J`�RR`jɽ�*<e�9����d����F��j(�d�A�ɽ�*<eɽ�*<e�ߐuX�q�-�]�x�r8��6ɽ�*<e��CQ�Ը�]_��;U�S�rh�ɽ�*<eg���Xd����F�����L��fVA�0 yɽ�*<e"�2ܡF��l-�^�� �q�����ɽ�*<e�7�_��E")��Ҝ�$(�dL	��D2�Fp�AA��'I�5ž Nb '�̖g�%���ɽ�*<e_:�>ŧ[��g�0�r6V/'>а�ɽ�*<e�׽��J�}=�;!���~�L���ɽ�*<e�+ �0��hQڱx��aiUj)��}ɽ�*<eɽ�*<e���t+Q�y/)��l;��Q�onv>�v2DaZqON9�-(�/�Ww���n&V�ɝ�����-�~�F���g�$���j�Tu?4��ي�`�4ji�t`��4r�Q�r�M�%�G��?"(�UKx2�֑]>��mI�z�#-K7�3]N|��r)d`b��\�()�Ľ.�Dz�.���U�ۄ��6n��=f�.��F{Kɽ�*<e�/���%󬱖����(8�|q{+�bt�A-�� 0��%rɽ�*<eɽ�*<e1? ��6�+t�c�K�]��s�kɽ�*<eɽ�*<eɽ�*<e����n��rɽ�*<e��ܑ��h"z<�'~�f7=.��ɽ�*<e�/���%���7�1��W���[�&�E�?9D�uǎqh��gn(`m�R#z�͌�?�(<���p�.��ͣj|�2�F6��j�/�-Ȳ�N�#ɽ�*<e[��ղ�fǇz��X3�v����W����
���2�h
�K=4ɽ�*<eY[v�_�ɽ�*<e5�?��
��;�d ��Hk�P��|�W����sp�ɽ�*<e��{Y\iqS��c�P ��E��6�J�EL�cm�m�����ɽ�*<eҝ[��R�ɽ�*<e�LOG۳=���f���2�a��/5��bhF_ɽ�*<eyh�S
cP��ry�k��堒�c����g�#wF��@�OG�ɽ�*<eNM{9q��ɽ�*<e�r�璉�.����>W�_�4�Gײ�,�IM�+�I���>Է4[��ղ�fǇz��X3�v����W�������h��UI��Iɽ�*<eY[v�_�ɽ�*<e�Gy6+�$�,�IM�+�IV�x�S����p��,ɽ�*<eX��~?�W#8�|q{+�?�{�/z����c��kQ�]�Q�Mɽ�*<e����n��rɽ�*<e+�n�/�G<��0�eg�/���b��M&ɽ�*<ex�r%=YF��)�xoĪ�K��ƐΝ����%�:ɽ�*<eɽ�*<e�����ɽ�*<e�����^��{fs��.v�f>;�݃����!��/���%�n�>�B"�kC����J��!㣝˻�%e�܉f��Iă�A�VJUT���?�(<��ɽ�*<e7[��İ��f�Ӗ�F>�w�LV�/�"�l��Z=�ɽ�*<e[��ղ�fǇz��X3�v����W��k|~.�pɽ�*<eɽ�*<eY[v�_�ɽ�*<e!�T9����#%N��R���7��$`љR�$����sb7��ɇ�F�$W.����|�.k-���!Eg2�����Q�]�Q�M,4���?wɽ�*<eɽ�*<e0��葠�Q���Д4��k���C��!I�2ɽ�*<ex�r%=YF��)�xoĪX�(��8
cJ_���Q�]�Q�Mɽ�*<e�����ɽ�*<e�]Ӟv�߷G�eyk���C�ɽ�*<eɽ�*<ex�r%=YF��)�xoĪX�(��8
c�"C�Ӏɽ�*<eɽ�*<e�����ɽ�*<e�]ӞvF��Պ�����<���^������Mh�Y��2�K+���H��6�Sd�~�fT��9��I��5�2-ɽ�*<ex�\�uɽ�*<e�X���4�Y���<���^��Y�Ű�\�kܥ��qɽ�*<e$����sb7��ɇ�F�$W.����|ZO��>t �ău�Y�'ɽ�*<e,4���?wɽ�*<eɽ�*<e���$�*�_Ҋo;�e�j�<�U�qɽ�*<eyh�S
cP��ry�k���~��!�AE
!�ɽ�*<eɽ�*<eNM{9q��ɽ�*<eH�*��h�A)���Im�Y��# N��ɽ�*<e$����sb7��ɇ�F�$W.����|uNK�[����h
�K=4ɽ�*<e,4���?wɽ�*<eɽ�*<e�#f̨�~ܚ�C����m�B���wo�	h�[��{Y\iqS��c�P����v�G5�td'�b�]���ɽ�*<eҝ[��R�ɽ�*<eg*D����Vm�B���V�D�VO]=Su���eɽ�*<e�����	�1�ϱ����bӶ��9�^8�7ɽ�*<eɽ�*<e����n��rɽ�*<e�N*z+N����`K�f�"���Nd"�O��ɽ�*<e=�i>�N�|80�2AVQPXp�P�Q�]�Q�Mɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��K��@�����s��Q�!I�2ɽ�*<e�����	�1�ϱ�1m e��\U�>:�ɽ�*<eɽ�*<e����n��rɽ�*<e+�n�/�G�߷G�eyf��}J!W-V8��+ Zɽ�*<eD�d�2u� ���ƙ"�#F��8����T�ɽ�*<eɽ�*<e�����ɽ�*<e8�q�ѱ�V8��+ Zu��Aı�i���<���^������Mh	�?�o�.��c��y�-۱�*�jCe�V8��+ Z�h
�K=4ɽ�*<ex�\�uɽ�*<e�m�v�����<���^7)�ĝfһ��K�`ɽ�*<ew�;L�::{���	���=pl?4��_jk�#��ɽ�*<eɽ�*<e,4���?wɽ�*<eɽ�*<e������_z+Q4�Q�I>/�4	(yaf��ٿ�Y��2�K+���H��6�Sd�~�fT^�0��şAwo��o�ău�Y�'x�\�uvS+ё@j�����T���Ş��i�5�MP��..+`��ɽ�*<ex�r%=YF��)�xoĪZm��B��H�@�p1�AE
!�ɽ�*<e�����ɽ�*<e�Ef�]��_z+Q4�QMlZp
T�m�B���dZ��`R�$���H��6�Sd�~�fT^�0��ş{M�y0��bm�B���*c�n��&ɽ�*<e"Rݗ]T��G5�td'�e#<�޼ů5�MP��˃�6��Rb�-�э�g�x�r%=YF��)�xoĪZm��B��H�@�p1˃�6��Rb��33��0�����ɽ�*<e�e	�5S�B���@%�q\+m"�GZ�V�sɽ�*<eyh�S
cP��ry�k��8�����w�=*~*���Vɽ�*<eNM{9q��ɽ�*<e���P��o����pÙEǛ'��d��-QJX��~?�W#8�|q{+�?�{�/z����P�V?�	��Щ/�Q�]�Q�M����n��r����2��"-ct賤`K�fnL����a+��c�ɽ�*<e��{Y\iqS��c�PZ�?�v&i5�m�3'k:��h��ɽ�*<eҝ[��R�ɽ�*<e��K��@��\�L{�������^EG5�td'���e0t8�|q{+�?�{�/z����P�V?� �^J��yϦM�|.{� ̛#ɽ�*<e+�n�/�G�����d<��pR0NnL����a����%�#��U��Z��{Y\iqS��c�PZ�?�v&i5~��/��K�am@��m�����ҝ[��R�ɽ�*<eP�ay��b���4�Qp?}&��׶�}SD+�?M�49�iv ([��ղ�fǇz��X3�ݥ D���z}x���Q�w�	�6�cɽ�*<eY[v�_�ɽ�*<e�������Ѧ�����X�Bh�W��.����A؊����]�찴�}0�@Z���ŗ AM��jtU��&�}�h
�K=4,4���?w����M�%Y�g�E����$�*?Ѳչ���7Ց�X2��~`��r\_*X�#~v'�w�֬���AV�n��NJ��� ..
A���ɽ�*<eNM{9q��ɽ�*<eH�*��h�AJ���$F��X�Bh�WC'�K��wȀ�3+����]�찴�}0�@Z���ŗ AM��jtR����m�Q�]�Q�M,4���?wɽ�*<eɽ�*<e�#f̨�~8l��	�%Y�g�E�D��ݹ�VdE�0(|�:B�2ƍ�zC�M�L�+���s$)�=�B $�ɽ�*<eҝ[��R�ɽ�*<ed��1�d.��H|��k=<R|=-4Wj̼�д������8�|q{+�?�{�/z�p�^(]e��C�]�Nf��h+�0�����n��r����M�d��j���ڳ�`K�f8l��	�L�����`..+`����{Y\iqS��c�P/��+�ͼ�f���9TI��~-y7�h
�K=4ҝ[��R�ɽ�*<e��K��@���>�dS@<R|=-}��&�rSX��~?�W#8�|q{+�?�{�/z�p�^(]e��A ��%�y���������n��rɽ�*<e+�n�/�G�߷G�ey���n��M^��i�?ɽ�*<e�����E-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e7��{��������ѩ���c�n_(VAߝ�c��.�$� Ӆ<§T��vU)�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT��ȅ5�+�!m>��e6�ڡ����Ve:�X��\��g�����6��n��_Lq f�&�������Y���:cl ��C��z󚅔��Q}���5�lcnNMG���뿓�؋��Ŵ�����e��Ċ�|�J���ɽ�*<e��pJ�1�7�A�7e���5�-��)ӕyƛ�R�n�8s6��ZL	��D2�.���)V��w�o傏(�Q3X,�+ �0��L��P�a��M�G�1�2Zs��Q,��.���)V�GT��)��S����{�+ �0��L��P�a��t�W����_����mQ��.���)V�yA�ߠ��j�;�y	�L�q�_�L��P�a�ĭ��l���v�����R���.���)V��|�������	z�i�j��lp���O��y�������H��6�Sd�~�fT��R(EC 0��%rɽ�*<e�/���%��8[����9(ύ��Bɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���MO�~Iy'p�k�ɽ�*<eX��~?�W#���N�^�gn(`m�R�lJ��j�<@�ͼ4���*l�����7F'�]h��p�.��ͣj|�2�Fz҄�����������X��~?�W#8�|q{+�?�{�/z����P�V?C{u�h��@ɽ�*<e����n��r����@��և�`��$�%�ܧ�	\�j�<�U�q�Y��2�K+���H��6�Sd�~�fT ��w����ᦲc�ɽ�*<ex�\�uɽ�*<e�m=����9�n��4�}j&��1�«Y��2�K+���H��6�Sd�~�fT ��w���Av�'�Bɽ�*<ex�\�uɽ�*<e���$�*K�K����̸B���"���w�N���H��6�Sd�~�fT ��w���"�#F��8����T�x�\�uɽ�*<e����o���S�B���@%yeTQ}��V8��+ Z�Y��2�K+���H��6�Sd�~�fT ��w����"vЅ\��b�]���x�\�uɽ�*<eن�\�)�e#<�޼ż�l�G��ɽ�*<eyh�S
cP��ry�k��8�����w�=*~*���Vɽ�*<eNM{9q��9�C�)���J�= ȉ>|
ϒ���ɽ�*<e��{Y\iqS��c�Paa24�2G7����ᦲc�ɽ�*<eҝ[��R��`���{�"M��
��U�����ɽ�*<e��{Y\iqS��c�Paa24�2G7���Av�'�Bɽ�*<eҝ[��R�!�T9�k����S櫼��'����V8��+ Z��{Y\iqS��c�Paa24�2G7���"�#F��8����T�ҝ[��R�"`�cd �!�(I켇y��k~�G������r#��U��Z��{Y\iqS��c�Paa24�2G7����"vЅ\��b�]���ҝ[��R���#)ϫ��K�am@������Ȣ���
���2�/���%���U�?��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���	D��:�^�����%����/�"�l��Z=ؓ��z:�-q26�\�ɽ�*<eɽ�*<eɽ�*<eɽ�*<ej	�%w\������~�W%8n��Y�f�.�ɽ�*<e(�B)�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eu;�Qݷ�2U���m)�[��/���?��a�磅"��Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곞�&`I��i`X�F��Ҩ��Y��/eJR�k�/eJR�k�/eJR�k�/eJR�k��h
�K=4)�,3u�A��e6�ڡJR�^���,>�1��O���a\!�����l�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�f�]&��,�l�~�«�u���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�����/�\U9��8P�,[h�
�+ɽ�*<eS�;��$�Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<e��M�R��Lc ����U�O'��U�A�/���%��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���	D��:�^�����%X2��(s��;QC�q�����z:�-q26�\�ɽ�*<eɽ�*<eɽ�*<eɽ�*<ej	�%w\�����TZm��I�
>zby"ɽ�*<e��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eu;�Qݷ�2U���m�|6*]�&��Jd�q/ݖ+ �0��MK�s�Zɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ��n�D2�B�"����ߛ	p�_�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ����Ve:�X��\��ݑ��/�׸s7��s�����Ɯ�h�[�Z�~�q��0��Y"�����Q��V��~�*.���HE")��Ҝ)*z�8$h�#��IJ<�+ �0���&9p��b8iS�0��)���m��M8����0E�\[$E")��ҜsN��8H��!���pXoXֺ��	w�F�#��ި}E](����Ðjɽ�*<embv��'0��]_��;.�w <>k��h����8�!�I*��d����F��#��V��~x !��ɽ�*<e�YA_٢`��T<�2�+�F��ɽ�*<eFiăU�?�E")��Ҝ��~�1�7��V��V��Fp�AA�A;��i���tgv
�i�S�DJɽ�*<e���㡆�.�, ����ჭ�u�lL	��D2)��O�WJh^ӽ6ԓ܌����c�9��-�/���%�����t\�M-�]�x�+� {�E�ɽ�*<e�X�C)�˸�]_��;�E�I6�H�T��qT�2y��d����F�6�_� �nɽ�*<eɽ�*<e�HA�?ݥG߬�:ǄA�>�M���!Tɽ�*<e?=���bZ2E")��Ҝ"CA��e���l�O�p�!:�{��@A;��i\�`�P�J�����G��Zɽ�*<e�/��{q�n9�F�c¾-L��vYmI�z�#-K��L���eEh^ӽ6���A��<�s��il��/���%�-�ٚ����3�Գ�fVA�0 yɽ�*<eٓ� �bѺ��jx���J��3"/��ɽ�*<e��U�ۄ��h^ӽ6Ԏm����kL	��D2�/���%��eG��Z-�]�x����g$�@ɽ�*<e8�Cc��S������\��;��+;�ɽ�*<e���뾚�d����F�����L�� �G?�L��ɽ�*<eʞ(�yh�=IG����u��]��ɽ�*<e�D�ů�ƟE")��Ҝ�$(�dH�T��q�Fp�AA��5D@/V���&�-����,	4ɽ�*<ek��1A���l�d�t������n�0�ɽ�*<e�0Q\��DU��b� ���1�p%�F�ɽ�*<e�+ �0��\�g?�.�3�	A��ŏ=����V��+ɽ�*<e���İ��z��｟��s���=u�^u��s�U��h��9ڡ�����@t����,�A�gҟVbw?,���L��P�a���ER�WV)���^Hɽ�*<e�ߐuX�q�g�M�9�mćX�V�?`�mI�z�#-K�.���)VA��F\���S�<v��%lɽ�*<eؕ�U�I�kDj��^��,Fwp�_c��x��'ѳ��w��ɽ�*<eɽ�*<e��+�J^�Q��	�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q��ɽ�*<e^��
:�*�~�sh-�ߠwo�	h�[ɽ�*<e�Y��2�K+��Qݓ˟s4�)�_π ����������'�e����Ǆ9�<7������r�<%:�=~<���%�6���s��Ɩ#�˴��56ɽ�*<ex�r%=YF�����?���D�	��}�o���ɽ�*<eɽ�*<e�����ɽ�*<e&O{��?=o��0Z������D�\å�)�}^Dz$����sbRIꐦO�j$W.����|Y�<d�2!#	76
m�"�ɽ�*<e,4���?wɽ�*<eɽ�*<e��"�m�+߀M:�`xr�a\� R�E���/���%�|2w�e�Q��kC�����ݮ5q.I<����<Q�]�Q�M�VJUT���?�(<��ɽ�*<e)_�6-�p�V�*��#E�����1��#�sɽ�*<ex�r%=YF�����?�ч�t}�,�IM�+�IQOB-�y�ɽ�*<e�����ɽ�*<e���|���(zSȢ�|N)�/Ԁ;�DhY��F�ɽ�*<eyh�S
cP�^��,Fwp�堒�c�!�}�>�ɽ�*<eɽ�*<eNM{9q��ɽ�*<eb4�j�d��gŬ/���?��ɽ�*<eX��~?�W#��	�d�?�{�/z�eg�/��y�����ɽ�*<e����n��rɽ�*<e+�n�/�G/���?��jKfz=��_d�Ǹ������-��Y��2�K+�I�\�m��`�f ��{�f>;�݃����h��Q�]�Q�Mx�\�uɽ�*<e�H��g澁_d�Ǹ��#��6*+�'��s<%��ɽ�*<eɽ�*<ex�r%=YF�����?�K��Ɛ��dsv��Zɽ�*<eɽ�*<e�����ɽ�*<e�bv�t>W�2Y��?ڼ%��9���wo�	h�[[��ղ�fǁ����=�v����W���R���7���՞WS�ɽ�*<eY[v�_�ɽ�*<eZi��LύE��9����;��i���!�)�49�iv (X��~?�W#��	�d�?�{�/z�k���C�w�	�6�cɽ�*<e����n��rɽ�*<e+�n�/�Gi���!�)�/V}�9�8mk��畬�ɽ�*<eX��~?�W#��	�d�?�{�/z�k���C��h
�K=4ɽ�*<e����n��rɽ�*<e+�n�/�Gl� �J��1Q����fٰ���˫�ɽ�*<e��{Y\iq���Lt�c�+[�&�����<���^��y���C�ɽ�*<eҝ[��R�ɽ�*<e��{��s����4�Qp?�*���U ��:��*�ɽ�*<e[��ղ�fǁ����=�JP�>��Av�'�Bɽ�*<eɽ�*<eY[v�_�ɽ�*<e!�T9���	3�Zq��()zӺ_gɽ�*<e�/���%�|2w�e�Q��kC����#E<[�hAf��Iă�Aɽ�*<e�VJUT���?�(<��ɽ�*<e��_NN��#3J�f)�������ɽ�*<e[��ղ�fǁ����=�JP�>���^ {�Eɽ�*<eɽ�*<eY[v�_�ɽ�*<e���������k_�:#_�"�#F��8#��U��Z$����sbRIꐦO�j$W.����|O\�;���m�B���m�����,4���?wɽ�*<eɽ�*<e����o���S�B���@%y�] �E�j&��1��ɽ�*<e�F`��� ^�k�Oڴf����.�NH�h
�K=4ɽ�*<eɽ�*<eNM{9q��ɽ�*<eX��zF��
��З�������P�ɽ�*<ew�;L�::{���	��v8��Z(8..
A���ɽ�*<eɽ�*<e,4���?wɽ�*<eɽ�*<e�m=����9M�(=��49�iv (ɽ�*<e�F`��� ^�k�Oڴf�ŏ�T��qQ�]�Q�Mɽ�*<eɽ�*<eNM{9q��ɽ�*<e���P���@!��dҠ����d<������of�����	�1�ϱ����~DB�!�(I���33��0ɽ�*<e����n��rɽ�*<e+�n�/�G�����d<��pR0N���U�'
Rٰ���˫�ɽ�*<e=�i>�N��utm&Y���v��{�5�2-ɽ�*<eɽ�*<eҝ[��R�ɽ�*<eP�ay��b���4�Qp?��'s��J�J=���ɽ�*<e�PI߬H����%hJT72�����j�D������ɽ�*<eɽ�*<eY[v�_�ɽ�*<e�2R&�N5݄p��P2��6�2��4\�kܥ��qɽ�*<e��{Y\iq���Lt�c�aa24�2G7���Av�'�Bɽ�*<eҝ[��R���j�Р��2�h	��`�\k�h}!�Lڜ�j�<�U�qX��~?�W#��	�d�?�{�/z���"o��D�$@�՛�f��Iă�A����n��rɽ�*<e+�n�/�G���q��6�2��4"�#F��8#��U��Z��{Y\iq���Lt�c�aa24�2G7���"�#F��8����T�ҝ[��R�ɽ�*<eg*D����Vm�B������}2�K��r�=_V8��+ ZX��~?�W#��	�d�?�{�/z���"o��D�Z�9�V8��+ Z�7F'�]hɽ�*<e+�n�/�G˃�6��Rbr�++�����^�s�H*��b��M&�/���%�|2w�e�Q��kC����m�@�-�F�^�� ���y������VJUT���?�(<��ɽ�*<e:��8*$7�He����ҟg'P��S(yaf��ٿyh�S
cP�^��,Fwpyyֶ�T@ÙEǛ'�h+�0�ɽ�*<eNM{9q���5��[1gԟ��R����HB����}x���Q�..+`��$����sbRIꐦO�j$W.����|�TErǃ++��c��h
�K=4,4���?wɽ�*<eɽ�*<e�m=����9He�����Z�j"�nm�B����Zc?Y��t^��,Fwpyyֶ�T@����^EG5�td'�b�]���NM{9q��ɽ�*<ew[i����Ç̸B����d=�#�<d}x���Q�˃�6��Rbsw�@�u!�RIꐦO�j$W.����|�TErǃ+����%�����T�,4���?wɽ�*<eɽ�*<eن�\�)�e#<�޼ń��P�V?�|L\h&�ɽ�*<ex�r%=YF�����?Ш6�E�SD+�?M��&ZReX�ɽ�*<e�����ɽ�*<e�� Qx����r=hJ��
ѥ䰾M^�������@�v;�z���v������D�Oȝ��QL�~PW:�=����ɽ�*<e�!4pL��X�Bh�W(�s:<�\��	3�Zq��[V�`���>Q����Ӆ<§Tg�����6��o�����:�X4 P��<1��M
�����VJUT���?�(<��ɽ�*<e��_NN���r=hJ��
ѥ䰾M^�^p�!P�@�v;�z���v������D�Oȝ��QL�~Pw�	�6�cɽ�*<eY[v�_�ɽ�*<e�������Ѧ�����X�Bh�WJ8�-�3!L7�Z^]��O]�찴�}0�@Z���ŗ|ptjy��zI�-�k��h
�K=4,4���?wɽ�*<eɽ�*<eM�Uy-V9?Ѳչ��&�����ڧ\�kܥ��qyh�S
cP�^��,Fwp���W�X��<R|=-4Wj̼��ău�Y�'�X�tJi��X�Bh�Ww=���`�O��lk��X�Bh�Wd��ٰ#s�����#i�RIꐦO�j$W.����|c� k�k��L�����`�AE
!�,4���?wɽ�*<eɽ�*<e�m=����9?Ѳչ��&�����ڧY��# N��yh�S
cP�^��,Fwp���W�X��<R|=-}��&�rS�h
�K=4NM{9q��ɽ�*<e���P��/V}�9�8\#����r�ɽ�*<e��d�r"�:Dx��pɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r���	$���2U���m5�:�]X��M��cD'�IYU��)�ٛR��@ZLK|�#ɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�u�
O]�S�7�V�B�f��+1��"��IpN��h�.�o��Ɗ�Iג$OJ�7��D����'-�rEJ�H���vN������έ�I�x6���_��=��O����Jb@���;7Pb䡑�9������/���%�73��<}$c~�L���L��+�
7�3]N|�<���	����	/���/���%󬧁��ȉ�iFj>· �Vn���3�
���Wϓg��eB��ڧ�q�-�m��Y��Mu �;Ϋ��rc�\��g?�V��w�
���Wϓ�YEG�_5��X��>�}b>�Jsg����ȉ�i1����κ�=�V��7�3]N|�9ܲ_�l�3uUrD쇝�
��ۧ���ȉ�in�(�˃׵O�g��.p(�qʱt�s��y����Lt�c�aa24�wM[��vg'ѳ��w��ɽ�*<eǋ'H)�@w����a���h
�K=4ɽ�*<eɽ�*<eɽ�*<ex�\�u���r�<,�����K�����]ɽ�*<e�,��T"���`χ�a$����^�M�"�ds��R��6G�2���-l	*vӈ����
%:�=~<���%�6��Aiq��%ɽ�*<eyh�S
cP�^��,Fwpyyֶ�T@E%��D�&�y�����ɽ�*<eNM{9q���&X�o��*C���w9:;\B��ɽ�*<e��{Y\iq���Lt�c�Z�?�v&i5�m�3'k:��h��ɽ�*<eҝ[��R��`���{A`@5�A�!d!p*�~�ɽ�*<e��{Y\iq���Lt�c�Z�?�v&i5�H�:���9�^8�7ɽ�*<eҝ[��R�!�T9��v��J�}���:��e
ٰ���˫���{Y\iq���Lt�c�Z�?�v&i5Pn���&���!�(I���33��0ҝ[��R�"`�cd �!�(I켰��}���J��tL:W������of��{Y\iq���Lt�c�Z�?�v&i5~��/��K�am@��m�����ҝ[��R���#)ϫ��K�am@� Nzw�Y��# N���/���%�|2w�e�Q��kC����m�@�-�F�^�� ���y������VJUT���?�(<��PD��7�	��̲�E6�..+`��$����sbRIꐦO�j$W.����|�o�K��o�zG����}��h��,4���?wɽ�*<e�Ef�]���̲�E6�Su���e$����sbRIꐦO�j$W.����|�o�K��o�G�e�2� ���9�^8�7,4���?wɽ�*<e��t5��;��̲�E6������d<��#�����RIꐦO�j$W.����|�o�K��o��������!�(I�G�;8�;�/ɽ�*<e8�q�ѱ�V8��+ Z��̲�E6�˃�6��Rbsw�@�u!�RIꐦO�j$W.����|�o�K��o����-���K�am@�Z<�}U�'�ɽ�*<e�e	�5S�B���@%�u��|���-Ȳ�N�#sAyA/��6����[ɽ�*<eɽ�*<eɽ�*<eɽ�*<ej	�%w\������~�W%8n�B�K*�]�ɽ�*<e(�B)�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eu;�Qݷ�2U���m)�[��mk��畬��+ �0��MK�s�Zɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곑f�[��!<�ɠ)�Fi=�Z ���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ��`���)6�LQ{D���b��M&ݭ�:nB�r/eJR�k�/eJR�k�/eJR�k�ec�*�S��ɽ�*<e��s��Q�V�B�f�]&��,�gj�T�1'�� oحɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�����/�\U9��8P�|�� ����!i�#%}ʔʵ�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��M�R��Lc �<gcp2��y�k">z���/���%�ȣleg�׿ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���	D��:�^�����%Z�SB~���'ZC��������ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<ej	�%w\�����R��kq6v�_��I���ɽ�*<e(�B)�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eu;�Qݷ�2U���m��̲�E6�}�-��%�a�磅"��Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ�ih�/�_R��X�����{��Q�h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ��|�KLǍ�M�U�帶[��%�w/����4�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�f��+1܃��.�?g��3nQ�t��Ϡ�Ab=��K�X}(�K�r��UY��q��JFV-O�;8W�f�W��*��'��/x���O�*����J��}�eC��8�xWfb��W�>ph^ӽ6��ӸP�[$��fE��Q�U�����W��"�e��l��^���Q8���M?��Z���ޓ>h^ӽ6��J��}�e��e6����/���%�s�@�uV��ި}E](�h�#��IJ<ɽ�*<esXӭ�(����Sy1��\t{Đ��-��!�G�z�2�=�d����F��Q�2k{�ȃ�?i\ɽ�*<e���<�J��O1��	��VZ uD�L	��D2D�҈q��E")��Ҝ��~�1�7P�lb�(��Fp�AA��kIR�cr�j�����٦%?zɽ�*<e{�����Z�.�, ����ჭ�u�lH�T��q)��O�WJh^ӽ6�%���Nbqz�d'uV��/���%���jm�1-�]�x�{ ���(5%ɽ�*<e�xz1EAʼ���⥦�MS�����ɽ�*<eȻsO� d����F��eif���ɽ�*<eɽ�*<eCk�naB�7iJ	�y�ֶÙ)ٔ:�OFD[7�Kͮ_E")��Ҝ#nZ~�n�W66��u7���N�S�<�x\�`�P�J�+�G.���}ɽ�*<eħ�����9�F�c.�E>2�<Uɽ�*<e&f�jJ�6h^ӽ6�Z�-��K#ɽ�*<e�/���%�h�����H��3�Գ� �G?�L��ɽ�*<e�.���)V���bX�Zr����9!ɽ�*<e��}2��h^ӽ6Ԏm����kH�T��q�/���%����qBl�e�>��9�B��K�ɽ�*<eT<�� ������\��F�+Sxɽ�*<e�pl�E{d����F�`�� �P1s�j݇�M�uɽ�*<e��dj^��=IG������á���ɽ�*<e����:r�sE")��ҜsK''oB�ɽ�*<e���m#P���<�)3=����)D����tx�E�Bxɽ�*<e1������6�=�����<�tx�E�Bxɽ�*<e�[���¸Q����JJ���;�X��d`���N��/���%�6rF
�E��8/�2!�ӣ��$n@�9pی��d��JęŎ�&��݆5�EB�v%��KZ��
���Wϓ��B�������	H�%1#�,�vL��U�ۄ���!���7�%\�j׸'��^H�/���%�u �;Ϋ�
*ȲX�mI�z�#-Kɽ�*<e�8����;K�Raz�kC������OL,4杖�#ڄɽ�*<e�/���%��8[����9(ύ��Bɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<��G�x9��FE�&I��}Kg��@հɽ�*<eɽ�*<emD�ْ�dh89QN��hz�;3��PY���F��
�W���[�&`�ժH���ҝ[��R�@d����і[.�[����;��w��\��ɽ�*<eX��~?�W#��Jnj��?�{�/z��s��Ɩ	�q��IX;ɽ�*<e����n��rɽ�*<e��J���Δm��ڙ�UZL�\A��˾�[(ɽ�*<e[��ղ�f�ڇ��C�v����W���D�\å�ᝄ�Dsɽ�*<eY[v�_�ɽ�*<e�c��,R#u��˾�[(jT��_���W��#T�&ꬶ�R�Y��2�K+��+ v��`�f ��{`xr�an�����1wɽ�*<ex�\�uɽ�*<eA��V	{�A�W��#T�l�(��7�ɕ?kV7�(T�F(��X��~?�W#��Jnj��?�{�/z�E������K��(Z�ɽ�*<e����n��rɽ�*<e+�n�/�Gɕ?kV7��w�H������{�\w6�ɽ�*<e�/���%�;K�Raz�kC����̾���ܔ7]��s�kɽ�*<e�VJUT���?�(<��ɽ�*<e	���j���FZ����<�ɠ)�Fɽ�*<eyh�S
cP�Ɖ�D��0L�堒�c�/���?���h
�K=4ɽ�*<eNM{9q��ɽ�*<e���U�&4�K����!*�A�������T�O�Nd"�O����{Y\iq��;�T2� ���_d�Ǹ��..
A���ɽ�*<eҝ[��R�ɽ�*<e��]/߷�W��T�O��C�_@�"�d�;�ɽ�*<eX��~?�W#��Jnj��?�{�/z�&�d}�=cUQ�]�Q�Mɽ�*<e����n��rɽ�*<e+�n�/�Gg��	� �E�&�ϔ���5�7��dhɽ�*<ex�r%=YF�n�Rd%�;~�)�D?R��9���m�����ɽ�*<e�����ɽ�*<eN�����K5�B�����S�b��i`X�F�ɽ�*<eyh�S
cP�Ɖ�D��0L�堒�c�i���!�)��&ZReX�ɽ�*<eNM{9q��ɽ�*<em�}�����OG}Db���S�b�ޔ'd����ɽ�*<eyh�S
cP�Ɖ�D��0L�堒�c�k;c���xɽ�*<eɽ�*<eNM{9q��ɽ�*<em�}����������"vЅ\��a�k|jZ�$����sbt���̌$W.����||P����J�yϦM�|.Q�]�Q�M,4���?wɽ�*<e�ub���ن�\�)�e#<�޼�(��ʸG�ɽ�*<eɽ�*<ex�r%=YF�n�Rd%�;�Y�<4~��9�^8�7ɽ�*<eɽ�*<e�����ɽ�*<e��t5��;�Hn��F�����-�ɽ�*<e�Y��2�K+��+ v���Sd�~�fT�	Qo��Q�]�Q�Mɽ�*<ex�\�uɽ�*<eW���P�#��6*+�'ն��@�f�ɽ�*<eɽ�*<ex�r%=YF�n�Rd%��:�W�Ӡ��\U�>:�ɽ�*<eɽ�*<e�����ɽ�*<e�� Qx����H�3���!�(I켔-�э�g�[��ղ�f�ڇ��C�JP�>��"�#F��8����T�ɽ�*<eY[v�_�ɽ�*<e"`�cd �!�(I���wv�&;���7dɽ�*<e�/���%�H'b6]��O0�|W:�=����ɽ�*<eɽ�*<e�VJUT���?�(<��:j���+�k\+��N��X9�/ח�q]�iʳ1ɽ�*<e�PI߬H����IÎ��X�Y6�M
����ɽ�*<eɽ�*<eY[v�_�ɽ�*<e�`���{G�鱚b�xa�׍hCɽ�*<e�/���%�H'b6]��O0�|w�	�6�cɽ�*<eɽ�*<e�VJUT���?�(<��ɽ�*<e:��8*$7��%��G�,��̸B���������Mh�F`��� ^!M��ch�L�PlC�V8��+ Z�h
�K=4ɽ�*<eNM{9q��ɽ�*<ew[i����Ç̸B���7)�ĝfһ�"vЅ\��a�k|jZ�w�;L�::{���	���L$�z�g����<���^��y���C�ɽ�*<e,4���?wɽ�*<eɽ�*<eن�\�)�e#<�޼��hc�V�G�c�тɽ�*<eD�d�2u���^�'��K�`�h
�K=4ɽ�*<eɽ�*<e�����ɽ�*<e�5ŀ�@$�h�<��ܪ�.����A��:��*�$����sbt���̌$W.����|�o�K��o�G�e�2� ���9�^8�7,4���?wɽ�*<e��*�M��嫑�$�*�q\+m"���~`��rɽ�*<eyh�S
cP�Ɖ�D��0L�8�����w�=*~XEߵW�,Q�]�Q�MNM{9q��ɽ�*<eH�*��h�A�c��J��K"U�8?1A��!�(I�sw�@�u!�t���̌$W.����|�o�K��o��������!�(I�G�;8�;�/ɽ�*<eɽ�*<e����o���S�B���@%�q\+m"�|M��t+c�����ofyh�S
cP�Ɖ�D��0L�8�����w�=*~�V��P ���5�2-NM{9q��ɽ�*<e����Ħ�
V8��+ Z�_z+Q4�Q�;�Y��##ɽ�*<e�Y��2�K+��+ v���Sd�~�fT^�0��ş��l�G���h
�K=4x�\�uɽ�*<e��Ԫ�N�Ml��+aC~ ��w���\�kܥ��q�/���%�;K�Raz�kC����K��H7�g'P��Său�Y�'�VJUT���?�(<����P�V?�6}����}&��׶�}��hƁ�,�j�<�U�q[��ղ�f�ڇ��C�ݥ D���z}x���Q��AE
!�ɽ�*<eY[v�_�ɽ�*<e�`���{R�5`�� ��w���"�#F��8�o���J|;K�Raz�kC����K��H7Z�j"�nm�B���(�ZZZ���?�(<��ɽ�*<eB��gJ��A���4�Qp?}&��׶�}��f�M�
V8��+ Z[��ղ�f�ڇ��C�ݥ D���z}x���Q�˃�6��Rb��33��0Y[v�_�ɽ�*<e��#)ϫ��K�am@����}2�K�E%��D�&��b��M&X��~?�W#��Jnj��?�{�/z����P�V?C{u�h��@ɽ�*<e����n��rɽ�*<e+�n�/�G�߷G�eyp�^(]e����j�M�Su���e�ɏu��7)��S�5��ȺTa�/"���S@�ࣨSɽ�*<e(�V�3~_ѥ䰾M^����")���}hc�f���9TI'�09k� �)���-B�*�v2}&�PZ�n.{{3VUv�b��ᦲc�ɽ�*<ex�\�uɽ�*<eW���P�#��6*+�'p�^(]e����j�M��!I�2�ɏu��7)��S�5��ȺTanW8����&ZReX�ɽ�*<e�����ɽ�*<e�� Qx����r=hJ��
ѥ䰾M^��i�����@�v;�z���v������D�Oȝ|�G�~�����u,ɽ�*<eY[v�_�ɽ�*<e�ܡ�,�'!I^�
��[V�`��,\�8� 'z,�ӻ��;K�Raz�kC����^��N2�{�&�����ڧAv�'�B�VJUT���qN4��T:TM�B"�O�@c��l2!�r=hJ��
TM�B"�Ol>j�m�[��ղ�f�ڇ��C������3e�X�Bh�Wd��ٰ#sf��Iă�AY[v�_�ɽ�*<e�`���{R�5`���[V�`���S�)n%�"C�;K�Raz�kC����^��N2�{�&�����ڧ�^ {�E�VJUT���?�(<��ɽ�*<e:��8*$7��WG��Kгj����N0ɽ�*<e8\(�U�M��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q����=�wYh�ǵ�r�k�7����f�y������&8_UXec��
ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�����/�\G�P�1�	��=#c?�V�Y��H�r��Ob��i���sX!�x���њJ'�R5�+ұ�"���k#�B�j�^9����CNh!�SM�oXֺ��	�2�����F�+��jd��)��\|}��i��K��ͳ[2�aEi7|2d>7L	��D2�ߐuX�q���#B����M�<h���U��h���Lw��Qv��J�ɽ�*<e}���5�lҐ��z��(]kM�U��h���qH �a���Ph��Bf���I�U�Z�}���5�lNӹqs�<$�l=�F���B�B�Lw��O0���O~,!�j��\�ߐuX�q�����Ph�n����ç^�^��^�Lw�群�	���xv.?���g�s�HB	�kt���̌$W.����|�o�K��o���N��-(���#ڄɽ�*<e��=!��(2��p�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�-��fΡ��k��4t�pԖ�����Mh�/���%���7�1��W���[�&�E�?9D�uǎqh��gn(`m�R#z�͌���od�t�[.�[����V���/��!I�2�/���%�;K�Raz�kC����K��H7E������h
�K=4�VJUT���?�(<�슂�s!貓�r�sc<5����-�$����sbt���̌$W.����|�TErǃ++��c��h
�K=4,4���?wɽ�*<e�Ef�]��zh#��d��-QJ$����sbt���̌$W.����|�TErǃ+�\�r+�=��h
�K=4,4���?wɽ�*<e��t5��;LӚٿr-�G5�td'� =��jB�t���̌$W.����|�TErǃ+3��|��V8��+ Z1wg�i"yPɽ�*<e8�q�ѱ�V8��+ Z��Moi��v���<���^185G��t���̌$W.����|�TErǃ+����%�����T�,4���?wɽ�*<e�e	�5S�B���@%o;���5���������Y��2�K+��+ v���Sd�~�fT^�0��ş��l�G���h
�K=4x�\�u]�P�.�F�#f̨�~?+�o&[��j�<�U�q[��ղ�f�ڇ��C�`E���փ<�~v3��>|
ϒ����h
�K=4Y[v�_�+�n�/�G���q���=X�Soj&��1��[��ղ�f�ڇ��C�`E���փ<�~v3����U������h
�K=4Y[v�_�+�n�/�G��`K�f��9üI`�̸B���'�UO���ڇ��C�`E���փ<�~v3�����'����V8��+ Z�iE����n+�n�/�G�����d<��pR0N� j�Y��V8��+ Z[��ղ�f�ڇ��C�`E���փ<�~v3��G������r����T�Y[v�_�+�n�/�G˃�6��Rb��wv�&ZP���t�o#�˴��56�f170
\Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<eu;�Qݷ�2U���m)�[��"�d�;��+ �0��MK�s�Zɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곞�&`I���'d������{��Q�h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ��`���)6�l���SI������������l�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�f|f��lW�^|��]`�g���X�mZ �/eJR�k�/eJR�k�/eJR�k�6����[����n��r�����/�\U9��8P�Y!���n ��S��v>�^1�?q�-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��M�R��Lc �Ij�a�*�QW+�_�����gY��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���	D��:�^�����%��jg�s��	�6���z:�-q26�\�ɽ�*<eɽ�*<eɽ�*<eɽ�*<ej	�%w\�����TZm��I�8K����ɽ�*<e��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eu;�Qݷ�2U���m��Moi��v��МB\'��+ �0��MK�s�Zɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ�\�)eE�;QC�q��i=�Z ���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ}X}�+5����K�`ɽ�*<e-&J�� ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�f��������Jd�q/ݏe��>� ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�����/�\G�P�1�	��=#c?��Z�ØKρ�XcQtp�)�پ������8B`}�FW,P���{Z��
�rt��l�-�b���~��4�1i�Jc2d����F��\	�je�1���b2ޏ� �G?�L��{ �L[�HzdI�4R��z��f��4.�����Sf�H���dd����F��A��~2��fҡ�^��L!�%��+�xՑ*�.�, ������b2ޏ�fVA�0 y�*����*"h^ӽ6��J��}�eC��8�xWf�/���%󬖡���2��
��
����f\�,�ɽ�*<e�u�;�"��]_��;��'g�;S1��<N]��q�����d����F����.ޛXSpL?l�ɽ�*<e�H�i3ﭠO1��	��VZ uD�H�T��q��qz�WE")��Ҝ�P��Ti��a
0�x�(�EqxP��E��ccr�j�����k�:?o
ɽ�*<e{�����Z����bX�ZH�c��ɽ�*<e��P�/�h^ӽ6�%���Nbq,1�Yބ��/���%�6� �����USm��]�fVA�0 yɽ�*<e�(	"<���⥦���G#��Cɽ�*<eT�-5F�nd����F��#��V�C�2w��Z[��!��bKٌ�٦7iJ	���y�j�(��aO�!��d�Տ�E")��Ҝ#"܇a��'~]����(�Eqx�j�Tu?4�\�`�P�J�ܒ��5H�ɽ�*<e[N����br�D�2;L	9��Fgɽ�*<e�
��Y�6�h^ӽ6�>�J#��(ɽ�*<e�/���%�j�Tu?4�:9y����B�p�?�ɽ�*<ex�g� ����bX�Z��A�a�l'ɽ�*<e[a�?~��h^ӽ6�Hk�K{�ԵL	��D2�/���%�j�$�'�Φe�>��9�̖g�%���ɽ�*<e���(�����jx���J���9��ɽ�*<ea�|xd����F�`�� �P1s��^!�]qɽ�*<e�jI�1�;ż��Q��R�k�!�ɽ�*<e��ލk�׫���;��ҟ�d	ɽ�*<es'Syo���<�)3=���K[�k�ɽ�*<eɽ�*<e/q���±�T�y:t�n�5Ǔ��G�tx�E�Bx%"	�E׋u:�`O;�~�T�ȭL���2�-g��H���gXF�+����꣺�X�#e<�P�XB�4M3}���5�l&2}��$sN��8H��ɽ�*<e�.���)VOL$���5�֎%;�#�,�vL�U��h��$�������a?���|\pɽ�*<e-��)ӕy��y�������]-��'5{��UĖZ�'[P�u�ɽ�*<eɽ�*<eǋ'H)�@w����a���h
�K=4ɽ�*<eɽ�*<eɽ�*<ex�\�uɽ�*<e�4����k���A�X:胮."1Do�ɽ�*<e$����sb����o=�����bC�x���b��6�-4�)�_πZ<�}U�'�:j���+�K�o��c�{��%B{$�"l�+���š�	"�$ɽ�*<eyh�S
cP�q>��Z�.�堒�c�)u/��L�<Q�]�Q�Mɽ�*<eNM{9q��ɽ�*<e	N�9���� 4���:o�QT�G!���s�-ɽ�*<ex�r%=YF�N'�����π�eפm���˾�[(�h
�K=4ɽ�*<e�����ɽ�*<e�Vz�+#} �h��x��[�y��aކ���jqɽ�*<e��{Y\iq��Ժ��h� ��E��6��W��#T�.�YСɽ�*<eҝ[��R�ɽ�*<e��&m�an����g�?�:p׌,㗟��<�Eɽ�*<eyh�S
cP�q>��Z�.�堒�c�ɕ?kV7�'~_�~Nɽ�*<eNM{9q��ɽ�*<eT��%��G㗟��<�E�4�ҷE��D�j�)Iɽ�*<e�Y��2�K+���]-��`�f ��{U���g(ɽ�*<eɽ�*<ex�\�uɽ�*<e?������ex���u�P�f>;�݃��������/���%󬖸3����kC����J��!㣝��v[o�I�^ɽ�*<e�VJUT���?�(<��ɽ�*<e7[��İ�����э�� ��P�6;7}�~�p[�3�$����sb�ϝO�}�$W.����|�z ��>���T�O�M
����,4���?wɽ�*<eɽ�*<eD���p �W"!��ٜ;��FZ����Nd"�O��ɽ�*<eyh�S
cP�q>��Z�.�堒�c�0ڧ�AO4ɽ�*<eɽ�*<eNM{9q��ɽ�*<e���U�&4��C�_@���rq��&�c���#�X��~?�W#|m9T�g�R?�{�/z��&�ϔ���2��Aqzɽ�*<e����n��rɽ�*<e+�n�/�G��rq��&�NB�q�vȮ�^q.J1��b��M&�/���%󬖸3����kC�����z��=D��M�N�ɽ�*<e�VJUT���?�(<��ɽ�*<e��DO�y4�{fs��.vr(HU�Qɽ�*<e�/���%󬖸3����kC�����z��=S�w��Rdɽ�*<e�VJUT���?�(<��ɽ�*<e�٣�eo��T#��Lg��K�am@��wo�	h�[[��ղ�f�������JP�>���"vЅ\��b�]���ɽ�*<eY[v�_�ɽ�*<e�E�$n�d�K�am@�c�ţ�`��Su���eɽ�*<eX��~?�W#|m9T�g�R?�{�/z�(��ʸG��h
�K=4ɽ�*<e����n��rɽ�*<e+�n�/�G��`K�f����qNd"�O��ɽ�*<e��{Y\iq��Ժ��h��LMǊ��..
A���ɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��K��@�BK�K�K�{�!I�2ɽ�*<eX��~?�W#|m9T�g�R?�{�/z�:�Y�e��Q�]�Q�Mɽ�*<e����n��rɽ�*<e+�n�/�G�߷G�eyw荦xy�cV8��+ Zɽ�*<ex�r%=YF�N'������6S�k�=�!�(I���33��0ɽ�*<e�����ɽ�*<e8�q�ѱ�V8��+ Zmm<�=T��d��-QJɽ�*<e	�?�o�.�z��d��Q.����T�3@�ࣨSɽ�*<eɽ�*<ex�\�uɽ�*<e�
�Ӛ�.����Ş��i9n��5�ɽ�*<eɽ�*<eD�d�2us��ĵ��&�ᦲc�ɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�Ef�]�'� ��h/��b��M&ɽ�*<e	�?�o�.�z��d��Q�0���Ѓ��&ZReX�ɽ�*<eɽ�*<ex�\�uɽ�*<e��Ԫ�N��iAfyl�ދF��ݕٰ���˫��/���%�H'b6]f2O]-Q�렽���d<��5�2-ɽ�*<e�VJUT���?�(<��ɽ�*<eB��gJ��A���4�Qp?0��l�-ǿ�K�am@��wo�	h�[�PI߬H��o,�)Nk��+��%�yϦM�|.Q�]�Q�Mɽ�*<eY[v�_�ɽ�*<e��#)ϫ��K�am@�V�D�VO]=,�o��vɽ�*<e�����	�1�ϱ�><���a.�"���ɽ�*<eɽ�*<e����n��rɽ�*<e+�n�/�G�ƚ�읶���]������ɽ�*<e[��ղ�f�������`E���փ<�~v3����U������h
�K=4Y[v�_�����2(�s:<�\��	3�Zq�B`�M����-��/���%󬖸3����kC����m�@�-�F�]��?�`C�..
A����VJUT���?�(<��ɽ�*<e��_NN�ζ���]�؊��SV8��+ Z[��ղ�f�������`E���փ<�~v3�����'����V8��+ Z�iE����nɽ�*<e"`�cd �!�(I�r�++�����/��Z �^���<���^[�Q��S���3����kC����m�@�-�F��I�|�ЮH���<���^#z�͌�?�(<��ɽ�*<eD$敃���pR0N6�2��4Y��# N��ɽ�*<e��{Y\iq��Ժ��h�aa24�2G7����^ {�Eɽ�*<eҝ[��R�ɽ�*<e�JLs�����_z+Q4�Q�H�:���:��*ȫY��2�K+���]-���Sd�~�fT ��w���Av�'�Bɽ�*<ex�\�uG�k`>-:���"��hρ��Ş��i���P�V?��a��{e�ɽ�*<ex�r%=YF�N'�����Ш6�E���hƁ�,f��Iă�Aɽ�*<e�����ɽ�*<e�Ef�]��_z+Q4�QPn���&���!�(I켥����TU���]-���Sd�~�fT ��w���"�#F��8����T�x�\�uɽ�*<e"Rݗ]T��G5�td'�e#<�޼ń��P�V?8����		%�����ofx�r%=YF�N'�����Ш6�E���f�M�
V8��+ Z�h
�K=4�����ɽ�*<e�e	�5S�B���@%He�����E�����ɽ�*<eyh�S
cP�q>��Z�.�yyֶ�T@E%��D�&�y�����ɽ�*<eNM{9q��ɽ�*<e���P��r"L�ń|%<R|=-�z�`u�tu1�D@u{�l�ʶ���u�[��|_�Nſ<�%K\�d�Q�]�Q�M����n��rp�^(]e���}��h����`K�f8l��	�%Y�g�E�����P�dE�0(|�:B�2ƍ�zC�ߕ�)��큰h��_�h��ɽ�*<eҝ[��R�ɽ�*<e��K��@���>�dS@<R|=-�n �u�HYaU�.n��p�l�ʶ���u�[��|_�Nſ2�1D���ɽ�*<e����n��rɽ�*<e+�n�/�G�߷G�eyp�^(]e����j�M�}�-��%��ɏu��7)��S��֧��`X�N�y��^C�U£���ɽ�*<e�����ɽ�*<e�����i���}hc�f���9TI���.�NH�Y��2�K+���]-���Sd�~�fT�[V�`��,\�8� 'z��9�^8�7x�\�up�^(]e��#ӛvn�J���Ş��ip�^(]e��#J�����`����-�x�r%=YF�N'�������㟰��TM�B"�OVQPXp�P�Q�]�Q�M�����ɽ�*<e�Ef�]����}hc�f���9TI�����7�Y��2�K+���]-���Sd�~�fT�[V�`���S�)n%�\U�>:�x�\�uɽ�*<e��Ԫ�N��{fs��.v2X0u0�pM*��U����/���%���U�?��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT��ȅ5�+�!m>��e6�ڡ�h�&u��p)2���@�h2uvÐ�2@�3�#[���HK
ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��p�^���Lc �v�l������4\���鳣���`��V�,�W]�ͻlU�� <�ZBg�cG4�NP�g���=z Ҡ�z;���ӷ�l2.��k���-F��lB��dzMp/�ar��\R`S�5�{AM�ɽ�*<e���[��c��#�����	/���U�ۄ���d���/)��H/��ɽ�*<ed��Ję���'�D&����A��tO�4�!���7�%�&�����V����Fd��Jęf5-�M0,�3��x�K���tO�4�!���7�%$�A��˼���d��Ję4��Wzhp�I�ۿww�佦i0Oh�!���7�%1�@ͫ�����e�ʝd��Jęs�Ϭ(�����Z){Q��r��<�-<���� �������`E���փ<�t�jA(OZ�'[P�u�ɽ�*<ew�;L�::=�Y��r����&6ɽ�*<eɽ�*<eɽ�*<e,4���?w:j���+�oaf�	��,��/�=X]ɽ�*<e�Y��2�K+��Qݓ˟s4�)�_π ����������'�e����ǄA�8���K�o��c�{��%B{$���}���49�iv (�Y��2�K+���]-���Sd�~�fT ��w���^ {�Eɽ�*<ex�\�u�&�|�D�#f̨�~a��#;�Nd"�O��[��ղ�f�������ݥ D���z}x���Q��AE
!�ɽ�*<eY[v�_�+�n�/�G���q��l2`�
��(yaf��ٿ[��ղ�f�������ݥ D���z}x���Q�W:�=����ɽ�*<eY[v�_�+�n�/�G��`K�f࣏�>�m�B���D���&�K������ݥ D���z}x���Q������d<��5�2-Y[v�_�+�n�/�G�����d<��pR0N���M���ٰ���˫�[��ղ�f�������ݥ D���z}x���Q�˃�6��Rb��33��0Y[v�_�+�n�/�G˃�6��Rb�y��k~�f��S�Hɽ�*<e��{Y\iq��Ժ��h�aa24�2G7����^ {�Eɽ�*<eҝ[��R�\/l�<�]��<}�l=2���mɽ�*<ex�r%=YF�N'�����Zm��B��H�@�p1�AE
!�ɽ�*<e�����H�*��h�Aa���d1�W�D6�fɽ�*<ex�r%=YF�N'�����Zm��B��H�@�p1W:�=����ɽ�*<e����옯��U�&4�h^�!�����ym��Aٰ���˫�x�r%=YF�N'�����Zm��B��H�@�p1�����d<��5�2-�����w[i����Ç̸B�����\>�_�V��P �޸����ofx�r%=YF�N'�����Zm��B��H�@�p1˃�6��Rb��33��0���������Ħ�
V8��+ Z)�[��w��\���:�<�.�ؙCB"��,#ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곑f�[��!Nd"�O����{��Q�h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ��`���)6�-�@v�ɽ�*<e-&J�� ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�f�б�͞8;7v��������pɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�����/�\U9��8P�6���N%��|�/��=1��[>�V�/eJR�k�/eJR�k�/eJR�k�,q'�Q�OQ�]�Q�M��M�R��Lc �Ij�a�*c�&�c���	����K��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���	D��:�^�����%��j��\�P�}7"\]e����,Wɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<ej	�%w\�����R��kq6v��%`���ɽ�*<e(�B)�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eu;�Qݷ�2U���m��̲�E6�y�k">z��a�磅"��Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곛�y�v|�iP��[P��{��Q�h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ��|�KLǍ�V����2ɽ�*<e�����l�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�f''�����J�J=���	���t�nj�'%萚 tɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�����/�\U9��8P�)�7h����X���W�
U�K;ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��M�R��Lc �v�l��Vh��S�zC��YB�gN2E[5���ԉ[��Q�)yӡ'�7�e�SuJg��/.�w <>k��h4�����#}w|�)�S�^5d�<l]j^a5k:e�."�v���l^��V���@}tV��^���>�A*��O2�9�L>2�kΟ���T�u�5�808;lAf ��)��v���l^�M��I�cr�j���[���K��ɽ�*<e)G;�?��I.�, ������b2ޏ� �G?�L����:Tǃ�h^ӽ6��IuW�������/���%�DY��x�v���f�9�O�����ɽ�*<e�jQK�6�	�y���:�S�Z�:���B�p�?� }�U�Pyd����F����.ޛ���1��ɽ�*<e�V/�P�R�p�Č�4�d���ɽ�*<e�Ewp��IE")��Ҝ�P��Ti��<��y�(�EqxP��E��c�"�YZR 6�q��ɽ�*<e��S�NW�ʵ��bX�ZE^�X,6�ɽ�*<e�Д��ʝh^ӽ6�Έ��"�q�ɽ�*<e�/���%��Y�Dxu��USm��]� �G?�L��ɽ�*<e1���\#����Sy1"�#$W&��L�0S0�?��<d����F��#��V�>Ey�U#�ɽ�*<e��$P/R�7iJ	��C�^a��ɽ�*<eyu��}��E")��Ҝu���|�����~M�D�(�Eqx�5D@/V��6�����L	��D2ɽ�*<e�;"���3r�D�2;LF�
('f�ɽ�*<e�U��h��E")��Ҝ � 	��#�ɽ�*<eL�@t�Z�s��V���@}:9y���}Mw�Ψɽ�*<e^iB�j�f��O�D d�4Oq��ɽ�*<e�k��)�h^ӽ6�Hk�K{�ԵH�T��q�/���%�S��\a�Z��p�q�xU�ީ�Lɽ�*<e� �;�m���jx���JMWK5�ޭ ɽ�*<ef�R�X6�Vd����F���'?�ڷI�tx�E�Bxɽ�*<e1M ҵ��[��^Us&�'2g�Doɽ�*<e%{5��0 ���Kx�?�^*���ɽ�*<e�v���l^N���Ir�nO9���c��LL�cɽ�*<e$Q0��0�{���`�)IjJ�+Rx��>�G�@7�3]N|��|���A��_�4��(���`�2]��tO�4�!���7�%fKˍʔ��	kU�f�Z�/���%󬧁��ȉ�id=MK(�b�sN��8H��ɽ�*<ed��Ję�� �2�ہ�-���ɽ�*<eY�9O=t�s��y�d��������~��]�H۝�ɽ�*<eɽ�*<e��=!��(2��p�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e�MO�~Iy'p�k�ɽ�*<eɽ�*<e[��ղ�f������ܛ�*l�����R��������sk��Y[v�_��K�{��e����F�5+!,D��(�q�
<~۞��>Է4�/���%���f�|L�kC����I�؊nޖ�,�\�ɽ�*<e�VJUT���?�(<��8�1���E��D�M�N�V�x�S���[�eonD+�'V��X��~?�W#;i���`C>?�{�/z��QT�G��J���:ɽ�*<e����n��rɽ�*<e+�n�/�G�[�eonD��gIU%٣�Д�٪,<Y��+�2$����sb(�2Y�ǫ$W.����|Fɱ�˕���2���}�ɽ�*<e,4���?wɽ�*<eɽ�*<eVd������ʴCj���>��܎��+dD�/���%���f�|L�kC�����Έx�3�㗟��<�E�h
�K=4�VJUT���?�(<��ɽ�*<e�|.���s��@B1}:��T��ɽ�*<eɽ�*<e��{Y\iqd������x���Y.w���`2���ɽ�*<eɽ�*<eҝ[��R�ɽ�*<eIh�����jKfz=�8;7v����ɽ�*<e�Y��2�K+�u�6�f�3`�f ��{�f>;�݃�\U�>:�ɽ�*<ex�\�uɽ�*<e�H��g澚c����w�LV�/���z�IYLy�q]�iʳ1[��ղ�fǕpᓖC�v����W���P�6;7}��]oT5��ɽ�*<eY[v�_�ɽ�*<e!�T9���z�IYLy�oc?3�<���4��6ɽ�*<e�/���%���f�|L�kC����J��!㣝�M
����ɽ�*<e�VJUT���?�(<��ɽ�*<e���,-a����� <�t-*�ɽ�*<eyh�S
cP�����N�B�堒�c���rq��&�������ɽ�*<eNM{9q��ɽ�*<e��{P���� <�t-*�5�:�]X^|��]`�ɽ�*<e�Y��2�K+�u�6�f�3`�f ��{Ȯ�^q.J1�y�����ɽ�*<ex�\�uɽ�*<e��vVK�`^|��]`�5�:�]Xf�af�w�ɽ�*<e�Y��2�K+�u�6�f�3`�f ��{˟M�o}Q�]�Q�Mɽ�*<ex�\�uɽ�*<e��vVK�`���;�	E��^��P#��U��Zɽ�*<ex�r%=YF����S,��m*?/�=Ȕ�K�am@��m�����ɽ�*<e�����ɽ�*<e'&���j�S�B���@%S�#�I.��j&��1��ɽ�*<eyh�S
cP�����N�B��~��!W:�=����ɽ�*<eɽ�*<eNM{9q��ɽ�*<e���U�&4�h��4��lR����P�ɽ�*<e$����sb(�2Y�ǫ$W.����|���t���M
����ɽ�*<e,4���?wɽ�*<eɽ�*<e�m=����9�Vt�� �g49�iv (ɽ�*<eyh�S
cP�����N�B��~��!w�	�6�cɽ�*<eɽ�*<eNM{9q��ɽ�*<e���P����g*l�<נ����d<������ofX��~?�W#;i���`C>?�{�/z�w荦xy�cV8��+ Z�h
�K=4����n��rɽ�*<e+�n�/�G�����d<��pR0N	6w���~w(yaf��ٿɽ�*<e=�i>�N��d�����IxL5�M�k/Q�]�Q�Mɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��Ӕh�75ÆJ|�㫘..+`��ɽ�*<e�����	�1�ϱ�4��U����h��ɽ�*<eɽ�*<e����n��rɽ�*<e+�n�/�G���q�����Y�B��ɽ�*<eɽ�*<e=�i>�N��d�����I2�ia�s�aɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e�JLs������+q)�;�G5�td'�a�k|jZ�	�?�o�.���k����W!`h FH�
�̸B�����y���C�ɽ�*<ex�\�uɽ�*<e"Rݗ]T��G5�td'�e#<�޼�O0�-x$�n#��U��Zɽ�*<eD�d�2u���ܠ�X��"vЅ\��b�]���ɽ�*<eɽ�*<e�����ɽ�*<e�e	�5S�B���@%fzA?���B�"���ɽ�*<e�F`��� ^�����ʽ��g�@P,͔�W�7�ɽ�*<eɽ�*<eNM{9q��ɽ�*<e$Ǟ�2ߊ$�l�	��p�5�MP��Su���eɽ�*<ex�r%=YF����S,��mZm��B��H�@�p1W:�=����ɽ�*<e�����<�B��Ѵ���")�_z+Q4�Q'�09k� �Nd"�O���Y��2�K+�u�6�f�3�Sd�~�fT^�0��ş91��?��M
����x�\�uɽ�*<eW���P�#��6*+�'�5�MP�⠽���d<������ofx�r%=YF����S,��mZm��B��H�@�p1�����d<��5�2-�����ɽ�*<e8�q�ѱ�V8��+ Z�_z+Q4�Q������^ٰ���˫�Y��2�K+�u�6�f�3�Sd�~�fT^�0��ştseQ,�yϦM�|.9�<7���ɽ�*<e�m�v�����<���^�d=�#�<dC'�K��wȶ������$����sb(�2Y�ǫ$W.����|�o�K��o���iMz�b�\U�>:�,4���?wɽ�*<eɽ�*<e�#f̨�~nL����a�\�r+�=�ɽ�*<e��{Y\iqd������Z�?�v&i5�H�:���9�^8�7ɽ�*<eҝ[��R���`�k�h���I6�{L�`�\k�h�����n������-�X��~?�W#;i���`C>?�{�/z����P�V?禺��zQ�]�Q�M����n��rɽ�*<e+�n�/�G���q��nL����a3��|��V8��+ Z��{Y\iqd������Z�?�v&i5Pn���&���!�(I���33��0ҝ[��R�ɽ�*<eg*D����Vm�B������}2�K��PO�K����<���^�%��Й�;i���`C>?�{�/z����P�V?8����		%�5�2-����n��rɽ�*<e+�n�/�G˃�6��Rbr�++���� ��w���Y��# N���/���%���f�|L�kC����K��H7E������h
�K=4�VJUT���?�(<��ɽ�*<e:��8*$7�?Ѳչ���7Ց�X2�ѥ����\_*X�#~v'�w�֬��n�r#�O1<�䴗�.�h+�0�ɽ�*<eN�����("<R|=-td������O��lk��X�Bh�W�	�y{I�7ع*i~x�h]�찴�}0�@Z���ŗZ������)�rj��+c�h
�K=4,4���?wɽ�*<eɽ�*<e�m=����9?Ѳչ���7Ց�X2GZ�V�s\_*X�#~v'�w�֬��n�r#�O1j�����0�y�����ɽ�*<eNM{9q��ɽ�*<e���P��r"L�ń|%<R|=-�;����ƃ�,�e��l�ʶ���u�[������/�P��!��Q�]�Q�M����n��rɽ�*<e+�n�/�G@ ^EZ�]8l��	�L�����`Su���e��{Y\iqd������/��+�ͼ�f���9TI���.�NH�h
�K=4��۩�f6<<R|=-��]2�f r�S�D�<R|=-��X�Y6������5C;i���`C>?�{�/z�p�^(]e��#J�����`..
A�������n��rɽ�*<e+�n�/�G���q��8l��	�L�����`�!I�2��{Y\iqd������/��+�ͼ�f���9TIŏ�T��qQ�]�Q�Mҝ[��R�ɽ�*<e�JLs����jKfz=��ڇ
�܎[ɽ�*<esAyA/��6����[ɽ�*<eɽ�*<eɽ�*<eɽ�*<ex�\�u�
O]�S�7�V�B�f���x4��Nl�>*�2�G���_D��{��QL�q�e���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_��MKZ�K������%C�k_�pw/�QL�L����A<NcM���N���Ɯ�h�[�Z�~�q�&��y�2�I����fRݵYi鸤(#�V�ƣ7�9<ځ8��$�z�ͺ}h���Z�dv�68�Fx�:�<�.�ص[1v��zyB=�u�@3M�<h���.���)V
��+���ŽA2�*PD-��)ӕyL��P�a���B���R��bT�>B�j�^9�V�U�M��$�L>d�-��)ӕy${t�|��h;��{f��.(�y/B�j�^9������71�y��i:,һ*�L��P�a�ē\[ ��J��4%~vD��.���)V��|�����j@��B���ǃ��lL��P�a�ĭ��l���vrR�\�\�k��=��h���Z0B�񇍞S,��mZm��B�]_+�w5�]�H۝�ɽ�*<e�
v�ƒm���X��cQ�]�Q�Mɽ�*<eɽ�*<eɽ�*<eY[v�_���ܑ��h"z<�'~�f7=.��ɽ�*<emD�ْ�dh89QN��hz�;3��PY���F��
�W���[�&`�ժH���a~va^�}l����F�P�T����)M E6N8Dɽ�*<e��{Y\iqd������Z�?�v&i5%�u�){K�\U�>:�ɽ�*<eҝ[��R�!��2����jN�̓������P�ɽ�*<ex�r%=YF����S,��mШ6�E���hƁ�,f��Iă�Aɽ�*<e�����H�*��h�A�5B�	��\�kܥ��qɽ�*<ex�r%=YF����S,��mШ6�E�.8��l@�ࣨSɽ�*<e����옯��U�&4�W�{�g��"�#F��8#��U��Zx�r%=YF����S,��mШ6�E��R�a�G��̸B�����y���C������w[i����Ç̸B�����,��"vЅ\��a�k|jZ�x�r%=YF����S,��mШ6�E���f�M�
V8��+ Z�h
�K=4���������Ħ�
V8��+ Z��̲�E6��!I�2$����sb(�2Y�ǫ$W.����|�o�K��o���iMz�b�\U�>:�,4���?w\Jԙ�% ��,���S!^����y�6����-�X��~?�W#;i���`C>?�{�/z���"o��D�$@�՛�f��Iă�A����n��rɽ�*<e��_NN���U�ݣ��d��-QJX��~?�W#;i���`C>?�{�/z���"o��D��Q(�>@�ࣨS����n��rɽ�*<e�0�i�X���,}�k�G5�td'���e0t;i���`C>?�{�/z���"o��D j��c�̸B���^0�\<efɽ�*<eB��gJ��A���4�Qp?��^� |����<���^�%��Й�;i���`C>?�{�/z���"o��D�Z�9�V8��+ Z�7F'�]hɽ�*<eD$敃���pR0N�D�pC���š�	"�$�>1�"@�q26�\�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ��`���)6C�b�MPɽ�*<e-&J�� ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�f|f��lW�f�af�w�	���t�nj�'%萚 tɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�����/�\U9��8P�F�.���!I�2�^1�?q�-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��M�R��Lc ��M��C!&���S+�"C��ʠ!4Nf/eJR�k�/eJR�k�/eJR�k��HTA��+�VJUT���	D��:�^�����%��j��\�J�����'��{
duzɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<ej	�%w\��������DC�MG�1G��ր͘�����A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eu;�Qݷ�2U���m��Moi��vΦ�-C��z�+ �0��MK�s�Zɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곮T.��͐�s��	�6i=�Z ���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ}X}�+5��D��ݹ�Vɽ�*<e-&J�� ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�f��^� |ҍ�МB\'�����pɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�����/�\U9��8P�ϰ1�d���G�c�тS�;��$�Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<e��M�R��Lc ����U�O��K�`�/���%�L�q�e���ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���	D��:�^�����%C�k_�pⳮ3f�d]HH��z�7DJq f�&�������E")��Ҝ)*z�8$���Ðj�+ �0���p'���:��0��Y"�����Q�����cn��ё�ǴJE")��ҜsN��8H��!���pXt�G��^*H�����b8iS�0��)���m7
s���H��%��+�{E")��Ҝ�����Q��V��~����m#P�͢j�Tu?4�cr�j���5k:e�."ɽ�*<ev��.�!9�F�c`ǌ����ɽ�*<e�����
h^ӽ6Ԋ6��_S�%���t�/���%�qAA|��!	�bđ;z��dI ɽ�*<e%�+�A�y���:�S�Z�:��}Mw�Ψ�S�|<1�d����F��� ����~��Ǡ/��^ɽ�*<e�Sñ8yYP�R�p�ČO𕓔��mɽ�*<e�Ewp��IE")��ҜΔ��B���fVA�0 y�(�Eqx�kIR��"�YZ/�ԂA�ɽ�*<e�r�:�N��螇�);D�ɽ�*<ep��T�5L`h^ӽ6Ԕ�j���3Kɽ�*<e�/���%�o�5�sc
��
���t�U�Y "�t��{d�.{�̎R����Sy1�CFG�؍N�}�*MO��As��ARFd����F��#��V�l�u?�u�ɽ�*<eo"�fxK��7iJ	�QC ��ӑɽ�*<e,��J>�jE")��Ҝ�˯.��ɽ�*<eL�@t�Z�s�5D@/V��6�����H�T��qɽ�*<ed��Ję.�n�	10c4�a�&r`ɽ�*<e޽\�4TE")��Ҝ����Njɽ�*<eL�@t�Z�sk�քM5�jv9��A��j݇�M�uɽ�*<e����|,�f��O�D���6sy�ɽ�*<e&0>����Sh^ӽ6�����H
��fVA�0 y�/���%�ڣ�	C�cQ��p�q�q�����ɽ�*<e�SX�:�������\�z}v�?�vɽ�*<e��K/�n^Tg��W���>R}9�ܲ��]iL�/���%󬎼�F��h���*b���]iLɽ�*<eI?��*��X�a���s�m]��ȋ��ϋ8z��L�@t�Z�sӟc�n��h|�%�9�m����k�ER$g#`��ߐuX�q��QF��V��:��k��wv��B�j�^9�T(�<7����*���s��[�U��h���Lw��c����^pl	kU�f�Z-��)ӕy9`��W�1�.Aҭ Uɽ�*<eɽ�*<es�HB	�k�
T����$W.����|̹尮l;�DhY��F�ɽ�*<ew�;L�::=�Y��r����&6ɽ�*<eɽ�*<eɽ�*<e,4���?wɽ�*<e���r�<,�����K�����]ɽ�*<eɽ�*<eO��'��P�n�/ͻ�:||hy�6"pUw�����I�� �p�����L���xr��<I}����hd�m��"�,w#ɽ�*<e�Y��2�K+I�b�H�`�f ��{�q�
<~�QOB-�y�ɽ�*<ex�\�uɽ�*<ek��+I JE��] �, �|��"m�w_�}�X"nɽ�*<eyh�S
cP��
��S�V�堒�c��[�eonDS2��Y5��ɽ�*<eNM{9q��ɽ�*<eM�J:xc>���T�JX[u�̏sLЭ�b\	y`�ɽ�*<e[��ղ�f�H���5�v����W��Д�٪,EWP���ɽ�*<eY[v�_�ɽ�*<eY�I����b\	y`��a�q� �l�Lj}��#�˴��56�Y��2�K+I�b�H�`�f ��{�>��܎�E#L�@���ɽ�*<ex�\�uɽ�*<e��Ԫ�N��Lj}����0Z����+�T���ɽ�*<e$����sb�
T����$W.����|���p�w��h
�K=4ɽ�*<e,4���?wɽ�*<eɽ�*<eU�Z�H� �*�A������!I�2ɽ�*<e��{Y\iq�f��2� ���c�H�hoM�Q�]�Q�Mɽ�*<eҝ[��R�ɽ�*<e��]/߷�W�߷G�eyeg�/�b2�M/��Jɽ�*<ex�r%=YF�2h�L�&�_�K��Ɛ·�z�IYLy�h��ɽ�*<e�����ɽ�*<e�����^�b2�M/��JjKfz=��Gܟ�ê.ɽ�*<e�Y��2�K+I�b�H�`�f ��{AQ�OsJɽ�*<eɽ�*<ex�\�uɽ�*<e�H��g�2$��Z�!�I����!�r칌,���/���%��/�ӄi�4�kC�������ʝ�u� <�t-*��h
�K=4�VJUT���?�(<��ɽ�*<e����{	b?�يq��r�k�7���|�/��=1ɽ�*<e��{Y\iq�f��L����^|��]`��h
�K=4ɽ�*<eҝ[��R�ɽ�*<e��r���
�JP$�r�k�7��&ꬶ�Rɽ�*<e��{Y\iq�f��L����!��pX��ɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��r�ϋ���WzM˃�6��Rb�-�э�g�X��~?�W#e���I?�{�/z���^��P����T�ɽ�*<e����n��rɽ�*<ec}��a�˃�6��Rbr�++����;���7dɽ�*<e�/���%��/�ӄi�4�kC����:���0r�=@�ࣨSɽ�*<e�VJUT���?�(<��ɽ�*<e�0�i�X󔑚�b�G�q]�iʳ1ɽ�*<e[��ղ�f�H���5�JP�>���ᦲc�ɽ�*<eɽ�*<eY[v�_�ɽ�*<e�`���{R�5`��xa�׍hCɽ�*<e�/���%��/�ӄi�4�kC������ޔ��	3�&ZReX�ɽ�*<e�VJUT���?�(<��ɽ�*<e:��8*$7��D#����̸B���������Mhyh�S
cP��
��S�V��~��!�����d<��5�2-ɽ�*<eNM{9q��ɽ�*<ew[i����Ç̸B���7)�ĝfһ\�kܥ��qɽ�*<ew�;L�::{���	��WWнm��h+�0�ɽ�*<eɽ�*<e,4���?wɽ�*<eiԙ�&�Vb���$�*~)�4hK���j�<�U�qɽ�*<e�F`��� ^�yC�~|5��~-y7�h
�K=4ɽ�*<eɽ�*<eNM{9q��ɽ�*<eH�*��h�A!���o��oY��# N��ɽ�*<ew�;L�::{���	���AY�����y�����ɽ�*<eɽ�*<e,4���?wɽ�*<eɽ�*<e�#f̨�~��G�=6m�B���wo�	h�[=�i>�N�Z�I�]�4j�s|Oݽ�yϦM�|.Q�]�Q�Mɽ�*<eҝ[��R�ɽ�*<eg*D����Vm�B���V�D�VO]=˃�6��Rb�-�э�g؟����	�1�ϱ�-f��`I��K�am@��m�����ɽ�*<e����n��rɽ�*<e+�n�/�G˃�6��Rb��wv�&�JzN̪[��%�w/�/���%�H'b6]{��S�~�o����7`Q�]�Q�Mɽ�*<e�VJUT���?�(<��ɽ�*<e�����E���/���z�`u�tj&��1��X��~?�W#e���I?�{�/z���"o��D��Q(�>@�ࣨS����n��rɽ�*<eA�G�]b�볤`K�f6�2��4����P�ɽ�*<e��{Y\iq�f��aa24�2G7����ᦲc�ɽ�*<eҝ[��R�ɽ�*<e��K��@��\�L{���c�XO�_ag�̸B���%��Й�e���I?�{�/z���"o��D j��c�̸B���^0�\<efɽ�*<e+�n�/�G�����d<��pR0N6�2��4�"vЅ\��a�k|jZ���{Y\iq�f��aa24�2G7����"vЅ\��b�]���ҝ[��R�ɽ�*<eP�ay��b���4�Qp?����]�^p�!Pɽ�*<e[��ղ�f�H���5�`E���փ<�~v3���t�s1�Q�]�Q�MY[v�_�ɽ�*<e��������N�Ky/�}x���Q�Su���e$����sb�
T����$W.����|�TErǃ+�\�r+�=��h
�K=4,4���?wvS+ё@ ��w��󃫑�$�*He�����Mc(J ��Nd"�O��yh�S
cP��
��S�Vyyֶ�T@�����n��..
A���ɽ�*<eNM{9q��ɽ�*<eH�*��h�A�c��J��K}x���Q������d<��#������
T����$W.����|�TErǃ+3��|��V8��+ Z1wg�i"yPɽ�*<eɽ�*<e����o���S�B���@%He������B5+o=�ٰ���˫�yh�S
cP��
��S�Vyyֶ�T@��PO�K����<���^��y���C�NM{9q��ɽ�*<e����Ħ�
V8��+ Z�_z+Q4�Q%�u�){K��������Y��2�K+I�b�H�Sd�~�fT ��w���^ {�Eɽ�*<ex�\�uɽ�*<e��Ԫ�N�Ml��+aC~�[V�`��G	�ģ�BH���N��g�����6��o����-V�P����d��2��.ău�Y�'�VJUT���Y�ǱE47�7Ց�X2���h��j��r=hJ��
ѥ䰾M^� b���@�v;�z���v������D�Oȝ2:(�@Հ�AE
!�ɽ�*<eY[v�_�ɽ�*<e�`���{R�5`���[V�`���>��h�
�$�:9���g�����6��o����-V�P�����))��h
�K=4�VJUT���?�(<��ɽ�*<e:��8*$7�?Ѳչ���7Ց�X2-�]K�T�*\_*X�#~v'�w�֬��2:���f~�{M)���Ǜ���ƑPiɽ�*<eNM{9q��ɽ�*<e4r�k�\���F���X�Bh�W.����T�3w�37+�
T����$W.����|c� k�k��L�����`W:�=����,4���?w{���0U_]&�����ڧ���$�*?Ѳչ��&�����ڧ����P�yh�S
cP��
��S�V���W�X��<R|=-��X�Y6�M
����NM{9q��ɽ�*<eH�*��h�AJ���$F��X�Bh�W�0���Ѓ�@%����g��
T����$W.����|c� k�k��L�����`w�	�6�c,4���?wɽ�*<eɽ�*<e�#f̨�~�h�������c�ޞ책ɽ�*<e�f170
\Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�����/�\U9��8P�k���C�\#����r�..+`��K��c��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e7��{���������R
�CI���$�$�w�'����ڎXNt���։Xb=��K�X}(�K�r��Z��T��U���Ɔ[E9錎��%�G��z�KZU���eh�V���v���l^���D8�*���xL	��D2^Gʵ��*�v1�g?�͸8yw�T��/���%�u �;Ϋ��}�{H����)��\|}�7�3]N|�T��@,j ��H"ԣ�|�/���%�o^H��(�B�7��~�$#rQ��ԚT7�3]N|������X���2��/���%�o^H��(�B_��-ϓG*u���7�3]N|�ڳ�f��-򲥎�w�-5�{�����ȉ�in�(�˃�5
I�S��Yk���E�9ܲ_�l �.�A�M[C�@��������(e���I?�{�/z���"o��D̹尮l;�DhY��F�ɽ�*<eg��1-P��V]��%�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����^��
:�*�~�sh-�ߠwo�	h�[$����sb����o=�����bC�x���b��6�-4�)�_πZ<�}U�'�L���xr��<I}�ԩ6�ֺ6��b��M&$����sb�
T����$W.����|�TErǃ+W=CՂ�z�Q�]�Q�M,4���?wɽ�*<e�w��ѹ����)��Y�q]�iʳ1X��~?�W#e���I?�{�/z����P�V?禺��zQ�]�Q�M����n��rɽ�*<e��_NN�΢jET�%���:��*�X��~?�W#e���I?�{�/z����P�V?�	��Щ/�Q�]�Q�M����n��rɽ�*<e�0�i�X�z�V���!�(I��^��j�e���I?�{�/z����P�V?� �^J��yϦM�|.{� ̛#ɽ�*<eB��gJ��A���4�Qp?��&�E@s��K�am@��m9C?'n�e���I?�{�/z����P�V?8����		%�5�2-����n��rɽ�*<eD$敃���pR0N�<�����49�iv ([��ղ�f�H���5�`E���փ<�~v3���t�s1�Q�]�Q�MY[v�_�^�����߷G�ey91��?��Nd"�O��yh�S
cP��
��S�V�8�����w�=*~XEߵW�,Q�]�Q�MNM{9q��W���P�#��6*+�'Awo��o�(yaf��ٿyh�S
cP��
��S�V�8�����w�=*~3�^�&��Q�]�Q�MNM{9q���H��g澁��Ş��i{M�y0��bm�B����Zc?Y��t�
��S�V�8�����w�=*~�ym��AyϦM�|.,K�%-
+["Rݗ]T��G5�td'�e#<�޼�tseQ,�ٰ���˫�yh�S
cP��
��S�V�8�����w�=*~�V��P ���5�2-NM{9q���m�v�����<���^�$ׁ��ݹE�=5�4���>Է4�����E-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�f�б�͞�Gܟ�ê.	���t�nj�'%萚 tɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�����/�\U9��8P�6���N%�&ꬶ�RS�;��$�Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<e��M�R��Lc ��M��C��P�6;7}2��S@�`��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���	D��:�^�����%e�2��B�$D�aSa>�p��Lf��/eJR�k�/eJR�k�/eJR�k�q26�\�j	�%w\��������DC�MX��Wo�������g��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eu;�Qݷ�2U���m�?ŸAl�Xȡ�m �G��y�Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ�f���t��(yaf��ٿ��{��Q�h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ��|�KLǍ+�����&ɽ�*<e�����l�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�f�S�{��%�u�d}l	���t�nj�'%萚 tɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�����/�\U9��8P��/1lG%iP��[P�^1�?q�-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��M�R��Lc �<gcp2��,�o��v�/���%�ȣleg�׿ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���	D��:�^�����%��`�l{�J�J=�������\	Mɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<ej	�%w\�����R
�CI���$�$�w�'�����j){��}��T��;.
�5�ג$OJ�7��D���O�*����J��}�e��e6���Xz2Y2�h^ӽ6���JFV-O�;8W�f��Y��M�]���%����l��^���Q8��;�#��l�,�yU�h^ӽ6��ӸP�[$��fE�ݾa8Z*�h��bo���s�P�R�p�ČO�;8W�fL	��D2 )�,.�E")��Ҝ�����Q�����cn��(�EqxA;��i\�`�P�J��wP��9�ɽ�*<eA�D�/?8�q���n`��r��E�
�*��@M�aɏ@xJ��h^ӽ6�J�k2����J��V2f�/���%��l�{R�F!	�bđxjt�ݯ�ɽ�*<eC�F���ƶ��]_��;�~�c�9hfVA�0 y �n8�]�d����F��� ����~��0�K��ɽ�*<e�Sñ8yY.�n�	10}o<]A�|�ɽ�*<e_�(/�Z�E")��ҜΔ��B��� �G?�L���(�Eqx�'I�5�øxQ@Q�;L	��D2ɽ�*<eӭ0��N����/'�6ɽ�*<eʡB��&yh^ӽ6�bN#D/Qi�W���8���}�i��{c���Ӫ
��
�������%ɽ�*<e{�O����B���Sy1o���R�-�	F��ݏ��������[d����F��#��V�>���u&D`ɽ�*<e��r�����{�h&��v@�.�1 ɽ�*<eB�Q�P�E")��Ҝ�Z��;���ɽ�*<e-��)ӕyd����F�{`is3Z�fVA�0 yɽ�*<ew�����s�.�n�	10�[m5t�ɽ�*<e-&�
:lݲE")��Ҝ��@��[�ɽ�*<e�Fp�AA��j�Tu?4�v9��A�􄘠^!�]qɽ�*<e�ˊ��'�?���n�0ilw|ɽ�*<eT6qRT*nh^ӽ6�����H
�� �G?�L���/���%󬦟�Ly�95�c�V壃.���|ɽ�*<e\�>ݺ-W��2�ٰj�!?�)�ɽ�*<e)����.g��W���P�.a7)�ɽ�*<e�/���%�q�>%��I��O�F��6���L�N�����]iL�I*{_���4{�〉6ᥘ2�
��0(�ڐ��U�ۄ���Z��x�yhɔ��|BjT;�9����(�C�x�o^H��(�BOD�ɕ�U�_rw���+ɽ�*<ed��Ję�,���,���=��Z���s��[7�3]N|���i�*��G�Y�ɽ�*<e��U�ۄ������ ��\�m0a��z��1�O'�;���ɽ�*<eɽ�*<e�
v�ƒm���X��cQ�]�Q�Mɽ�*<eɽ�*<eɽ�*<eY[v�_�ɽ�*<e-��fΡ��k��4t�pԖ�����Mhɽ�*<eX��~?�W#���N�^�gn(`m�R�lJ��j�<@�ͼ4���*l�����7F'�]h�G�x9��F�`둺��r�H9�����3�OZl(T�F(��ɽ�*<e��{Y\iq*��ř%(qS"�3�l�\[5���d�ɽ�*<eɽ�*<eҝ[��R�ɽ�*<e�~D�Uj�w�H�����A�c���ƁQu=�U��/���%���?��B��kC�����o�2��vc6%8�s���Q�]�Q�M�VJUT���?�(<��ɽ�*<e�Nl��h�Z/1�Q�W�wM�.����y֜�V���ɽ�*<ex�r%=YF����V���5�d��X,��b\	y`��h
�K=4ɽ�*<e�����ɽ�*<e��L��	�P�]��c�����U�:���y��Vɽ�*<e��{Y\iq*��ř%(94���i�Lj}��	�q��IX;ɽ�*<eҝ[��R�ɽ�*<e�t�<=��BDw��?p�����=/ʛ�_�wɽ�*<e[��ղ�f��\�m0a�v����W�����S�ɽ�*<eɽ�*<eY[v�_�ɽ�*<e�v�l�W]b]�
S4��P�6;7}49�iv ($����sb�s7�}��$W.����|�z ��>�w�	�6�cɽ�*<e,4���?wɽ�*<eɽ�*<eD���p �W/V}�9�8/���?��..+`��X��~?�W#�`���$��?�{�/z�eg�/�b2�M/��J�h
�K=4����n��rɽ�*<e+�n�/�G/���?�����q��*�A�����ɽ�*<eɽ�*<e��{Y\iq*��ř%(2� ���TD�>蔽iɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��]/߷�W5�:�]XM�L>�;>cW1	tqtV�Y��2�K+;	��7�8`�f ��{I����!����$e6ɽ�*<ex�\�uɽ�*<e��vVK�`M�L>�;>c�g�	>q�_!&���S+�������$����sb�s7�}��$W.����|̃��h�&,�v�1�V�ɽ�*<e,4���?wɽ�*<eɽ�*<e�4ł��滛�э�� �&�ӂ[uɽ�*<e$����sb�s7�}��$W.����|̃��h�&,.�YСɽ�*<e,4���?wɽ�*<eɽ�*<e�����I��rH�&V8��+ Zɽ�*<eyh�S
cP�r)1�ڹ���~��!˃�6��Rb��33��0ɽ�*<eNM{9q��ɽ�*<en�+E2�'V8��+ Z�8��.��ɏd��-QJɽ�*<e�Y��2�K+;	��7�8�Sd�~�fT�a��tO��Q�]�Q�Mɽ�*<ex�\�uɽ�*<e�H��g澁��Ş��iv�7�w�ɽ�*<eɽ�*<ex�r%=YF����V��؏��K���$�h��ɽ�*<eɽ�*<e�����ɽ�*<e�Ef�]�����Pk��b��M&ɽ�*<e�Y��2�K+;	��7�8�Sd�~�fT~��`��ɽ�*<eɽ�*<ex�\�uɽ�*<e��Ԫ�N�Ml��+aC~ދF��ݕٰ���˫��/���%���?��B��kC�����&u̿1�̸B�����y���C��VJUT���?�(<��ɽ�*<eB��gJ��A���4�Qp?�m����H��:��*�ɽ�*<e�PI߬H���q �y�4Wj̼��ău�Y�'ɽ�*<eɽ�*<eY[v�_�ɽ�*<ev�5�S;�{*�r�Ŝ�ÿ()zӺ_gɽ�*<e�/���%�H'b6]�)mh�%��AE
!�ɽ�*<eɽ�*<e�VJUT���?�(<��ɽ�*<e��_NN�Π��<�$V��������ɽ�*<e�PI߬H���q �y�}��&�rS�h
�K=4ɽ�*<eɽ�*<eY[v�_�ɽ�*<e���������f�fQI �"�#F��8#��U��Zw�;L�::{���	��5�%��č�G5�td'�b�]���ɽ�*<e,4���?wɽ�*<eɽ�*<e����o���S�B���@%]�)��x�V8��+ Zɽ�*<e�F`��� ^\ѯ
��?���W�������T�ɽ�*<eɽ�*<eNM{9q��ɽ�*<e����Ħ�
V8��+ Zk��� E����Jd�q/�ɽ�*<e	�?�o�.���R>W�G�i�.�!/O�|�*��ɽ�*<eɽ�*<ex�\�uɽ�*<e�ҋ\�d��6��V^��q\+m"��ѥ����ɽ�*<eyh�S
cP�r)1�ڹ��8�����w�=*~3�^�&��Q�]�Q�MNM{9q��G�k`>-:td������HB�����	�y{I�7�q]�iʳ1$����sb�s7�}��$W.����|�o�K��o�zG����}��h��,4���?wɽ�*<eɽ�*<e�m=����9�q\+m"��s��<��Gٰ���˫�yh�S
cP�r)1�ڹ��8�����w�=*~�ym��AyϦM�|.,K�%-
+[ɽ�*<ew[i����Ç̸B����d=�#�<d�J7�����K�am@��T��Fi��s7�}��$W.����|�o�K��o����-���K�am@�Z<�}U�'�ɽ�*<eɽ�*<eن�\�)�e#<�޼ů5�MP���!I�2ɽ�*<ex�r%=YF����V���Zm��B��H�@�p1w�	�6�cɽ�*<e�����ɽ�*<e�� Qx���}&��׶�}.8��lj&��1��[��ղ�f��\�m0a�ݥ D���z}x���Q�W:�=����ɽ�*<eY[v�_���j�Р���aH�M7u��	3�Zq� ��w�������P��/���%���?��B��kC����K��H7Mc(J ��M
�����VJUT���?�(<��ɽ�*<e��_NN��}&��׶�}�R�a�G��̸B���'�UO����\�m0a�ݥ D���z}x���Q������d<��5�2-Y[v�_�ɽ�*<e"`�cd �!�(I�r�++���� ��w����"vЅ\�J3�W�`>+��?��B��kC����K��H7�B5+o=�yϦM�|.��ZXd�"?�(<��ɽ�*<eD$敃���pR0NnL����a^ţ�U�ɽ�*<e��{Y\iq*��ř%(Z�?�v&i5%�u�){K�\U�>:�ɽ�*<eҝ[��R�ɽ�*<e�JLs�������}hc�f���9TI�I>/�4	HAD�j+��v2}&�PZ�n.{{��;���Av�'�Bɽ�*<erL۪w�Ib�[V�`��J�\4�^Ɂ��Ş��ip�^(]e����j�M�..+`���ɏu��7)��S����w�̈́���f�f��Iă�Aɽ�*<e�����ɽ�*<e�Ef�]����}hc�f���9TI�;�Y��##�m<>�m�^�v2}&�PZ�n.{{��;����^ {�Eɽ�*<ex�\�uɽ�*<e��Ԫ�N�Ml��+aC~�[V�`�����@��=�$�⥴F�1g�����6��o����f�c��O4����U�b9v�B	��VJUT���?�(<��ɽ�*<e&9��? �r=hJ��
TM�B"�O0��� �[��ղ�f��\�m0a������3e�X�Bh�W.����T�3@�ࣨSW�w:{&؁[V�`���SӜ�W\��	3�Zq��[V�`��zǙ�7�4Wu�?X�g��?��B��kC����^��N2�{�&�����ڧ�ᦲc��VJUT���?�(<��ɽ�*<e��_NN���r=hJ��
TM�B"�OE��4�[��ղ�f��\�m0a������3e�X�Bh�W�0���Ѓ��&ZReX�Y[v�_�ɽ�*<e�������Ѫ��э�� ������&ꬶ�R�:�<�.�ؙCB"��,#ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��p�^���Lc ��ӗEڔ����(�-����)P�hx#1w3mL��
�9�Հ�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r���	$���2U���m�  ƿzp�b�m���b�Ɏ���dF՘yӬ����8B`}�FW,P��=�����^O���	�%��.h�s�޼<����K!�R�Ժ����.f�_z�×��OK|��Qڨf���xɽ�*<e��x�>R}9�ܽA2�*PD�U��h���C�� $��0��<��f�ɽ�*<e�ߐuX�q�C��?�'�P�*�p'ݵYi��Lw��6UQ��/l��ܼ@"�ߐuX�q�u�:5jy��� �|I�tݵYi��Lw���`{����Be��	Qz�ߐuX�q�����w쑣�gW�Yi�p��~�@�Lw�群Ә��Aw�}�š/��ߐuX�q�����Ph=��t��oGs���9=I�kDj��r)1�ڹ��8�����꭭>���;���ɽ�*<e1? ��6�+t�c�K�]��s�kɽ�*<eɽ�*<eɽ�*<e����n��r�G�x9��FE�&I��}Kg��@հɽ�*<e[��ղ�f������ܛ�*l�����R��������sk����ss2�)��`둺��r�H9�����`�2�ɽ�*<e[��ղ�f��\�m0a�ݥ D���z}x���Q�w�	�6�cɽ�*<eY[v�_�)��6��l�߷G�ey�M`.�ɽ�*<eyh�S
cP�r)1�ڹ�yyֶ�T@�����n��..
A���ɽ�*<eNM{9q��W���P�#��6*+�'�F�W����ɽ�*<eyh�S
cP�r)1�ڹ�yyֶ�T@ÙEǛ'�h+�0�ɽ�*<eNM{9q���H��g澁��Ş��i�(���V8��+ Zyh�S
cP�r)1�ڹ�yyֶ�T@����^EG5�td'�b�]���NM{9q��"Rݗ]T��G5�td'�e#<�޼����q�ޤ#��U��Zyh�S
cP�r)1�ڹ�yyֶ�T@��PO�K����<���^��y���C�NM{9q���m�v�����<���^��\>�_��7zN-ɽ�*<ex�r%=YF����V���Zm��B��H�@�p1w�	�6�cɽ�*<e�����D��N_��^[V�Cg�����P��/���%���?��B��kC����m�@�-�F�]��?�`C�..
A����VJUT���?�(<���K��@��@��\�kܥ��q�/���%���?��B��kC����m�@�-�F��9�:~���h+�0��VJUT���?�(<����]/߷�W6�v����"�#F��8�o���J|��?��B��kC����m�@�-�F�4�)�*�z�G5�td'��C�	�?�(<��g*D����Vm�B��� Nzw��"vЅ\�J3�W�`>+��?��B��kC����m�@�-�F��I�|�ЮH���<���^#z�͌�?�(<��P�ay��b���4�Qp?3�w7]�'m��"�,w#��d�r"�:Dx��pɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�����/�\U9��8P�F�.��ɽ�*<eS�;��$�Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<e��M�R��Lc ��M��C�&�ӂ[u�/���%�ȣleg�׿ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���	D��:�^�����%����/�5�'��,������ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<ej	�%w\������~�W%8n��Y�f�.��!I�2gː�Ï��/eJR�k�/eJR�k�/eJR�k̩�o�w
H�ɽ�*<eu;�Qݷ�2U���m�?ŸAl�6Zg��7��~�,�~Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ�n���k��d���^���Ǘ����X��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ}X}�+5��'��U�Aɽ�*<e-&J�� ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�f��^� |�Φ�-C��z����pɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�����/�\U9��8P�y�C3-j4ɽ�*<eS�;��$�Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<e��M�R��Lc ����U�OD��ݹ�V�/���%��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���	D��:�^�����%e!ߖ�r�B�"������z:�-q26�\�ɽ�*<eɽ�*<eɽ�*<eɽ�*<ej	�%w\�����TZm��I�1�o%���G�c�тb��x���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eu;�Qݷ�2U���m�  ƿzp��'a�y�鍕D�3�/j�u�x��b��i���sX!�摠Z����\	�je�1���b2ޏ�fVA�0 yH�5��P�{Z��
�rt��l�-Z���Kza ׺{G��2d����F��A��~2��fҡ�^���%w��v�ߣ��}إ"zdI�4R��z��f��4.� *=5[0�Y�j�9Dd����F����:^���b���~��ɽ�*<e+���\�P�R�p�ČO�;8W�fH�T��qKV��G��E")��Ҝ����2�1��Eݤ/�(�Eqxk�քM5�j�:K�i��t���J}E�ɽ�*<e�l�Y�m��"�  v�C �7�fVA�0 y��xO&��h^ӽ6�J�k2����lg�f'%�/���%������H�ި}E](��^�����ɽ�*<eC�`�� ��]_��;�~�c�9h �G?�L�� �n8�]�d����F����:94�Pz��2��ɽ�*<e%���b`
_.�n�	10]�pTWɽ�*<e�:|�l��eE")��Ҝ�=�_�OU�ɽ�*<eu7���NP��E��cøxQ@Q�;H�T��qɽ�*<e������2�9�F�c����������撗wA�f��h^ӽ6�`q��Z�@T�R��n�/���%�@!!���
��
���-S��N�	ɽ�*<e����:�ـ��Sy1��T'ig���aO�!�M$�mVed����F�}D�4iɽ�*<eɽ�*<e��R�/�x{�h&��vP�5wu��ɽ�*<e7�3]N|���]_��;��Ox�nQ&ɽ�*<e.��x�y�Nd����F�{`is3Z� �G?�L��ɽ�*<e�A����חl-�^�� �xU�ީ�Lɽ�*<e�1q6�\
E")��ҜY;������ɽ�*<e���m#P��P��E��c� Nb '�B��K�ɽ�*<e���Pz%w�?���n���@� �ɽ�*<e��mp�n�h^ӽ6ԥ~3?7`����]iL�/���%�pP3�am���hAU6]?���,	4ɽ�*<e�#wƇv���C�g�{��tr��ɽ�*<e/�WA�Y0�{��NȈ�^�hq>Q��a�l��ɽ�*<e�%������En�]H��Q1���LHH0��.���)V�0�z���m��h{��6.b���ݵYi��Lw�羈�g���.�Dz�.�-��)ӕyL��P�a��$���$t�_rw���+ɽ�*<e�ߐuX�q�oL�P{�Pw\!h��m\ɽ�*<erP/�ۻ���Z0B��>���+�5K��#�����Xv�kɽ�*<eɽ�*<eg��1-P��V]��%�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�����:j���+�oaf�	��,��/�=X]ɽ�*<eɽ�*<e�,��T"���`χ�a$����^�M�"�ds��R��6G�2���-l	*vNM{9q����;��R�˴qZ5�����9u���
���2ɽ�*<e$����sbdf!п�$W.����|txG�z��h'~_�~Nɽ�*<e,4���?wɽ�*<e�Ja�f�ل�%�>v;�jT��_��J�EL�cm�wo�	h�[�Y��2�K+@w�����`�f ��{�A�c��ԃߔ�B���ɽ�*<ex�\�uɽ�*<eA��V	{�AJ�EL�cm��;�����g�#w�'�S 5l�X��~?�W#m��3+� �?�{�/z�wM�.�����$�c>y�Dɽ�*<e����n��rɽ�*<e+�n�/�G���g�#ww@&T.�f������h���+n��$����sbdf!п�$W.����|�� �"y&�sn5&;�Q�]�Q�M,4���?wɽ�*<eɽ�*<e���#B? ��T�i��6s��}�ɽ�*<eɽ�*<ex�r%=YF�>���+�5��8�z4ؓ���+4�ɽ�*<eɽ�*<e�����ɽ�*<e�h�z��qc�w�LV�/�5�'��,��ɽ�*<e[��ղ�f� �D�O�h>v����W���P�6;7}�&ZReX�ɽ�*<eY[v�_�ɽ�*<e!�T9�u�P�+H�"��FZ���ͻ�%e�܉�j�<�U�qyh�S
cP�C�6�vm��堒�c�/���?���AE
!�ɽ�*<eNM{9q��ɽ�*<e���U�&4��%e�܉�0����P��IPd��Qɽ�*<e$����sbdf!п�$W.����|�z ��>��h
�K=4ɽ�*<e,4���?wɽ�*<eɽ�*<eM��u�^8:㋞f����(H��u�6�ɽ�*<e��{Y\iq(�&��L����M�L>�;>cc��R��Mbɽ�*<eҝ[��R�ɽ�*<e�H�خ���v蛍::���x4��B�$Dɽ�*<e[��ղ�f� �D�O�h>v����W�!&���S+�\U�>:�ɽ�*<eY[v�_�ɽ�*<eșQ�z�~���;=6
����x4���QWk�HZ�ɽ�*<e[��ղ�f� �D�O�h>v����W�"���y��ɽ�*<eɽ�*<eY[v�_�ɽ�*<eșQ�z�~�к���@��9��I������of�/���%��x�#αh�kC�����<-`__�V8��+ Z�h
�K=4�VJUT���?�(<��vS+ё@�v�D�,��pR0N����Y�(yaf��ٿɽ�*<e��{Y\iq(�&���#ڴ-P�h+�0�ɽ�*<eɽ�*<eҝ[��R�ɽ�*<e��]/߷�W����G"l..+`��ɽ�*<eX��~?�W#m��3+� �?�{�/z�v�7�w��h
�K=4ɽ�*<e����n��rɽ�*<e+�n�/�G���q���&�M���ɽ�*<eɽ�*<e��{Y\iq(�&���,�)7�1��y�����ɽ�*<eɽ�*<eҝ[��R�ɽ�*<e�JLs����
�Y�7f�OG5�td'�a�k|jZ��Y��2�K+@w������Sd�~�fTދF��ݕyϦM�|.Q�]�Q�Mx�\�uɽ�*<e"Rݗ]T��G5�td'�e#<�޼�s$w�h�'ɽ�*<eɽ�*<eD�d�2u�� �O�Av�'�Bɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e��eZ�L�G��b�`�Ҧ���-�ɽ�*<e	�?�o�.�{.6���d��ٰ#sf��Iă�Aɽ�*<eɽ�*<ex�\�uɽ�*<eW���P�#��6*+�'n�E-��bɽ�*<eɽ�*<eD�d�2u�� �Oड^ {�Eɽ�*<eɽ�*<eɽ�*<e�����ɽ�*<e�� Qx��ӂ�c�H���!�(I켔-�э�g؀PI߬H��9�5P,�Ȍ���\�m�B���m�����ɽ�*<eY[v�_�ɽ�*<e"`�cd �!�(I���wv�&��9��I������of�/���%�H'b6];�\����˃�6��Rb��33��0ɽ�*<e�VJUT���?�(<��ɽ�*<eD$敃���pR0N���ᇴM��X���ɽ�*<e=�i>�N��6�$?��[���MĞ��ڭ�oqE�ɽ�*<eɽ�*<eҝ[��R�ɽ�*<e
�'63��ׇ�f���@
���B��d��-QJ�/���%��x�#αh�kC����m�@�-�F��9�:~���h+�0��VJUT���?�(<��^�u������h��j�����]� b��ɽ�*<e[��ղ�f� �D�O�h>`E���փ<�~v3��>|
ϒ����h
�K=4Y[v�_�ɽ�*<e�`���{R�5`�����P2��G5�td'J3�W�`>+�x�#αh�kC����m�@�-�F�4�)�*�z�G5�td'��C�	�?�(<��ɽ�*<eB��gJ��A���4�Qp?����]6vZ�%�M#��U��Z[��ղ�f� �D�O�h>`E���փ<�~v3��G������r����T�Y[v�_�ɽ�*<e��#)ϫ��K�am@����}2�K�n �u�HY49�iv (X��~?�W#m��3+� �?�{�/z���"o��D�2nq�Ř��&ZReX�����n��rɽ�*<e+�n�/�G�߷G�ey���P�V?TO�Ɩ�tzɽ�*<ex�r%=YF�>���+�5Ш6�E�.8��l@�ࣨSɽ�*<e������B֊ ��f�̚νEn�_z+Q4�Q�m�3'k:��q]�iʳ1�Y��2�K+@w������Sd�~�fT ��w����ᦲc�ɽ�*<ex�\�uɽ�*<eW���P�#��6*+�'���P�V?� �^J��ٰ���˫�x�r%=YF�>���+�5Ш6�E��R�a�G��̸B�����y���C������ɽ�*<e8�q�ѱ�V8��+ Z�_z+Q4�Q~��/��K�am@�dZ��`R�$@w������Sd�~�fT ��w����"vЅ\��b�]���x�\�uɽ�*<e�m�v�����<���^�d=�#�<d}x���Q��!I�2$����sbdf!п�$W.����|�TErǃ+W=CՂ�z�Q�]�Q�M,4���?wɽ�*<eɽ�*<e�#f̨�~8l��	�%Y�g�E�\�kܥ��qdE�0(|�:B�2ƍ�zC>��@��8�$�ss]d��9�^8�7ɽ�*<e�	��l\�f���9TI2�h	�r�S�D�<R|=-}!�Lڜh�8FP�G�l�ʶ���u�[����_��;��v믜�LQ�]�Q�M����n��rɽ�*<e+�n�/�G���q��8l��	�%Y�g�E�Y��# N��dE�0(|�:B�2ƍ�zC>��@��8�8�����}�\U�>:�ɽ�*<eҝ[��R�ɽ�*<e�JLs�������}hc�f���9TI�&!�r8�E�7��Ala�v2}&�PZ�n.{{�t�3�2���<�wj@�ɽ�*<ex�\�uɽ�*<e�m�v����>Ѷe%Ap�^(]e��C�]�Nf�ݏd��-QJx�r%=YF�>���+�5��㟰��TM�B"�OxL5�M�k/Q�]�Q�M��fT�u|f���9TI�9�k��˅��}hc�f���9TI��~-y7�Y��2�K+@w������Sd�~�fT�[V�`��zǙ�7��h��x�\�uɽ�*<eW���P�#��6*+�'p�^(]e��A ��%��b��M&x�r%=YF�>���+�5��㟰��TM�B"�O2�ia�s�aɽ�*<e�����ɽ�*<e�� Qx��ӵw�LV�/�u���vQ�jɽ�*<e�>1�"@�q26�\�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eY[v�_��MKZ�K������%��S�b��L{���V݅Ϗm�/
S�;��$�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q����=�wY�@o��W������&�5�D���z���'呝]A���C��&���Q�)y����-���F�ud�^jN�z/32�
���Wϓ���cp��RJlJ���ܡVx��a�l�/��/�8�0qe��]��c=���DХ�Oq�c�]�h�,�B��)��\|}�d��Ję���.���L��+�
��U�ۄ���!���7�%� Q��5ɽ�*<e�%�G��o�d�BjZ@L�cs���U�ۄ�����K�u�	H /�)w$[��ڱ��%�G����A�I�򄷘x������C�I��!���7�%0_S�do5���d��Jęs�Ϭ(�����C�K�e��	�!���7�%1�@ͫ����5)"�0��8�����x�#αh�kC����m�@�-�F�&�U �H����Xv�kɽ�*<e��+�J^�Q��	�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q���4����k���A�X:胮."1Do�ɽ�*<eO��'��P�n�/ͻ�:||hy�6"pUw�����I�� �pQ��/�%×�˴qZ5���,�Y��# N��ɽ�*<ex�r%=YF�>���+�5Ш6�E�SD+�?M��&ZReX�ɽ�*<e�����㵫�*�	�Z|[s%�o..+`���/���%��x�#αh�kC����K��H7Mc(J ��M
�����VJUT���?�(<���K��@�G5��3iv�Su���e�/���%��x�#αh�kC����K��H7�g'P��Său�Y�'�VJUT���?�(<����]/߷�W�LG�������d<�- �Ƈ����x�#αh�kC����K��H7Z�j"�nm�B���(�ZZZ���?�(<��g*D����Vm�B�����V���/�˃�6��Rb9k/�i����x�#αh�kC����K��H7�B5+o=�yϦM�|.��ZXd�"?�(<��P�ay��b���4�Qp?wb۳.��:��b��M&X��~?�W#m��3+� �?�{�/z���"o��D�2nq�Ř��&ZReX�����n��r���&B��G��θ��x�H�q]�iʳ1�Y��2�K+@w������Sd�~�fT^�0��ş91��?��M
����x�\�uɽ�*<e�m=����9í�>0\͟�:��*ȫY��2�K+@w������Sd�~�fT^�0��şAwo��o�ău�Y�'x�\�uɽ�*<e���$�*��́��>��!�(I켥����TU@w������Sd�~�fT^�0��ş{M�y0��bm�B���*c�n��&ɽ�*<e����o���S�B���@%;�� ����K�am@�dZ��`R�$@w������Sd�~�fT^�0��ştseQ,�yϦM�|.9�<7���ɽ�*<eن�\�)�e#<�޼ŝ� �v��(T�F(��8\(�U�M��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��M�R��Lc ��M��C�IPd��Q�/���%�ȣleg�׿ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���	D��:�^�����%e�2���QWk�HZܓ��z:�-q26�\�ɽ�*<eɽ�*<eɽ�*<eɽ�*<ej	�%w\������~�W%8n�Y��]��J��b��M&��A^ٿqɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eu;�Qݷ�2U���m)�[��i���!�)�!���rv�J3�tM/eJR�k�/eJR�k�/eJR�k�_�p�fh+�,4���?w��=�wYh�ǵ�n���k��d.e�&�ͮ�7��fc�Pɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡJR�^��hX�Wk�k�s����Od�����l�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�f?�
��#&'ZC��	���t�nj�'%萚 tɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�����/�\U9��8P�ɉj�]�!�(yaf��ٿ�^1�?q�-ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��M�R��Lc �<gcp2��}�-��%��/���%�ȣleg�׿ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���	D��:�^�����%����AYe�u�d}l������ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<ej	�%w\�����R��kq6vc���ġ[��%�w/(�B)�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eu;�Qݷ�2U���m��̲�E6�,�o��va�磅"��ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wY�@o��W������&�5G���0��Jf�x�\("��	�wR"]�ͻlU�� <�ZBg)�S�^5d�<l]j^a[���K���v���l^P��E��cSuJg��/.�w <>k��h����8��G�T�u�5�808;l>��J$�~�v���l^�'I�5�tV��^���>�A*�Ӭ��g0��@�D�b��]_��;.�w <>k��h4���5<�����d����F����:^��Z���Kzaɽ�*<e�?is���ئ7iJ	��qz�v�;ɽ�*<e=���5|+E")��Ҝ�}�9��F�Q�)(�Vx���m#P�͓�V���@}���tgv
�!#�Bw�ɽ�*<e�h����"�  v�C �7� �G?�L��zG��.�h^ӽ6ԓ܌���/%X@�S%�/���%�����t\�M�ި}E](�N��ɽ�*<eC�`�� ��]_��;�E�I6�L	��D2d��8���d����F����:94gإ���٣ɽ�*<e���a��N߬�:ǄA�hǳ�o�ɽ�*<e�]��Q��E")��Ҝ:���RTɽ�*<eL�@t�Z�s�kIR�\�`�P�J��b~*R�R�zr��A�lԃ��G�w9�F�c@�8�!5�/�w�Yݿ��h^ӽ6Զ�����֋R��D���/���%��.����G�
��
�����$S�ƾɽ�*<e�\�]�#����jx���J`�RR`jɽ�*<e�9����d����F��j(�d�A�ɽ�*<eɽ�*<e�ߐuX�q�-�]�x�r8��6ɽ�*<e��CQ�Ը�]_��;U�S�rh�ɽ�*<eg���Xd����F�����L��fVA�0 yɽ�*<e"�2ܡF��l-�^�� �q�����ɽ�*<e�7�_��E")��Ҝ�$(�dL	��D2�Fp�AA��'I�5ž Nb '�̖g�%���ɽ�*<e_:�>ŧ[��g�0�r6V/'>а�ɽ�*<e�׽��J�}=�;!���~�L���ɽ�*<e�+ �0��hQڱx��aiUj)��}ɽ�*<eɽ�*<e���t+Q�y/)��l;��Q�onv>�v2DaZqON9�-(�/�Ww���n&V�ɝ�����-�~�F���g�$���j�Tu?4��ي�`�4ji�t`��4r�Q�r�M�%�G��?"(�UKx2�֑]>��mI�z�#-K7�3]N|��r)d`b��\�()�Ľ.�Dz�.���U�ۄ��6n��=f�.��F{Kɽ�*<e�/���%󬱖����(E)�dC��z��1�O'�;���ɽ�*<eɽ�*<e�
v�ƒm���X��cQ�]�Q�Mɽ�*<eɽ�*<eɽ�*<eҝ[��R�ɽ�*<e�MO�~Iy'p�k�ɽ�*<eɽ�*<e[��ղ�f������ܛ�*l�����R��������sk��ҝ[��R�@d����і[.�[����;��w��\��ɽ�*<eX��~?�W#E)�dC��v����W����
���2�h
�K=4ɽ�*<eY[v�_�ɽ�*<e5�?��
��;�d ��Hk�P��|�W����sp�ɽ�*<e1��zfA�kC�����o�2��vc6%8�s���Q�]�Q�M�VJUT���?�(<��ɽ�*<e�Nl��h�Z/1�Q�W�wM�.����y֜�V���ɽ�*<ev���y�1�$W.����|Fɱ�˕���2���}�ɽ�*<e,4���?wɽ�*<eɽ�*<eVd������ʴCj���>��܎��+dD�/���%�c�i�#J?�{�/z�E������K��(Z�ɽ�*<e����n��rɽ�*<e+�n�/�Gɕ?kV7��w�H������{�\w6�ɽ�*<e�/���%�c�i�#J?�{�/z����c��kQ�]�Q�Mɽ�*<e����n��rɽ�*<e+�n�/�G<��0�eg�/���b��M&ɽ�*<ev���y�1�$W.����|�z ��>�w�	�6�cɽ�*<e,4���?wɽ�*<eɽ�*<eD���p �W/V}�9�8/���?��..+`��X��~?�W#E)�dC��v����W���P�6;7}��]oT5��ɽ�*<eY[v�_�ɽ�*<e!�T9���z�IYLy�oc?3�<���4��6ɽ�*<e�/���%�c�i�#J?�{�/z�&�d}�=cUQ�]�Q�Mɽ�*<e����n��rɽ�*<e+�n�/�Gg��	� �E�&�ϔ���5�7��dhɽ�*<ev���y�1�$W.����|�.k-���!Eg2�����Q�]�Q�M,4���?wɽ�*<eɽ�*<e0��葠�Q���Д4��k���C��!I�2ɽ�*<ev���y�1�$W.����|̃��h�&,�v�1�V�ɽ�*<e,4���?wɽ�*<eɽ�*<e�4ł��滛�э�� �&�ӂ[uɽ�*<e$����sbT��82�9`�f ��{˟M�o}Q�]�Q�Mɽ�*<ex�\�uɽ�*<e��vVK�`���;�	E��^��P#��U��Zɽ�*<ev���y�1�$W.����||P����J�yϦM�|.Q�]�Q�M,4���?wɽ�*<e�ub���ن�\�)�e#<�޼�(��ʸG�ɽ�*<eɽ�*<ev���y�1�$W.����|ZO��>t �ău�Y�'ɽ�*<e,4���?wɽ�*<eɽ�*<e���$�*�_Ҋo;�e�j�<�U�qɽ�*<e�+�
�na���g�_���K���$�h��ɽ�*<eɽ�*<e�����ɽ�*<e�Ef�]�����Pk��b��M&ɽ�*<e�Y��2�K+׷�����0��~��!w�	�6�cɽ�*<eɽ�*<eNM{9q��ɽ�*<e���P����g*l�<נ����d<������ofX��~?�W#E)�dC��JP�>��"�#F��8����T�ɽ�*<eY[v�_�ɽ�*<e"`�cd �!�(I���wv�&;���7dɽ�*<e�/���%�H'b6]2V���r�W:�=����ɽ�*<eɽ�*<e����n��rɽ�*<e�N*z+N����`K�f�"���Nd"�O��ɽ�*<e=�i>�N�Vnl�@�2�VQPXp�P�Q�]�Q�Mɽ�*<e�VJUT���?�(<��ɽ�*<e��_NN�Π��<�$V��������ɽ�*<e�PI߬H��n!B�dYo}��&�rS�h
�K=4ɽ�*<eɽ�*<eҝ[��R�ɽ�*<e�JLs������+q)�;�G5�td'�a�k|jZ�	�?�o�.��#���v!`h FH�
�̸B�����y���C�ɽ�*<eNM{9q��ɽ�*<ew[i����Ç̸B���7)�ĝfһ�"vЅ\��a�k|jZ�w�;L�::{���	���s*���|���<���^��y���C�ɽ�*<ex�\�uɽ�*<e�m�v�����<���^7)�ĝfһ��K�`ɽ�*<ew�;L�::{���	���n[�l��s�_jk�#��ɽ�*<eɽ�*<ex�\�uɽ�*<e�ҋ\�d��6��V^��q\+m"��ѥ����ɽ�*<e�+�
�na���g�_Zm��B��H�@�p1W:�=����ɽ�*<e�����<�B��Ѵ���")�_z+Q4�Q'�09k� �Nd"�O���Y��2�K+׷�����0�8�����w�=*~XEߵW�,Q�]�Q�MNM{9q��ɽ�*<eH�*��h�A�c��J��K"U�8?1A��!�(I�sw�@�u!�T��82�9�Sd�~�fT^�0��ş{M�y0��bm�B���*c�n��&ɽ�*<e"Rݗ]T��G5�td'�e#<�޼ů5�MP��˃�6��Rb�-�э�g�v���y�1�$W.����|�o�K��o����-���K�am@�Z<�}U�'�ɽ�*<eɽ�*<eن�\�)�e#<�޼ů5�MP���!I�2ɽ�*<ev���y�1�$W.����|�o�K��o���iMz�b�\U�>:�,4���?wɽ�*<eɽ�*<e�#f̨�~nL����a�\�r+�=�ɽ�*<e1��zfA�kC����K��H7�g'P��Său�Y�'�VJUT���?�(<����P�V?�6}����}&��׶�}��hƁ�,�j�<�U�q[��ղ�f���;��Y�Z�?�v&i5�m�3'k:��h��ɽ�*<eҝ[��R�ɽ�*<e��K��@��\�L{�������^EG5�td'���e0tE)�dC��ݥ D���z}x���Q������d<��5�2-Y[v�_�ɽ�*<e"`�cd �!�(I�r�++���� ��w����"vЅ\�J3�W�`>+�c�i�#J?�{�/z����P�V?8����		%�5�2-����n��rɽ�*<e+�n�/�G˃�6��Rbr�++���� ��w���Y��# N���/���%�c�i�#J?�{�/z����P�V?C{u�h��@ɽ�*<e����n��rɽ�*<e+�n�/�G�߷G�eyp�^(]e����j�M�Su���e�ɏu��7)��S��H!��/"���S@�ࣨS,4���?w����M�%Y�g�E����$�*?Ѳչ���7Ց�X2��~`��r\_*X�#~v'�w�֬�Ț�/�� ��NJ��� ..
A���ɽ�*<e�����ɽ�*<e�Ef�]����}hc�f���9TI�;�Y��##�m<>�m�^�v2}&�PZ�n.{{8�/���[�^ {�Eɽ�*<eNM{9q��ɽ�*<e���P��r"L�ń|%<R|=-�;����ƃ�,�e��l�ʶ���u�[����֙2Lx�P��!��Q�]�Q�MY[v�_�ɽ�*<e�ܡ�,�'!I^�
��[V�`��,\�8� 'z,�ӻ��c�i�#J?�{�/z�p�^(]e��C�]�Nf��h+�0�����n��r����M�d��j���ڳ�`K�f8l��	�L�����`..+`��1��zfA�kC����^��N2�{�&�����ڧ�ᦲc��VJUT���?�(<��ɽ�*<e��_NN���r=hJ��
TM�B"�OE��4�[��ղ�f���;��Y�/��+�ͼ�f���9TIŏ�T��qQ�]�Q�Mҝ[��R�ɽ�*<e�JLs����jKfz=��ڇ
�܎[ɽ�*<esAyA/��6����[ɽ�*<eɽ�*<eɽ�*<eɽ�*<eNM{9q����=�wYh�ǵ�r�k�7����f�y������&8_UXec��
ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT��ȅ5�+�!m>��e6�ڡ����Ve:�X��\��g�����6��n��_Lq f�&�������Y���:cl ��C��z󚅔��Q}���5�lcnNMG���뿓�؋��Ŵ�����e��Ċ�|�J���ɽ�*<e��pJ�1�7�A�7e���5�-��)ӕyƛ�R�n�8s6��ZL	��D2�.���)V��w�o傏(�Q3X,�+ �0��L��P�a��M�G�1�2Zs��Q,��.���)V�GT��)��S����{�+ �0��L��P�a��t�W����_����mQ��.���)V�yA�ߠ��j�;�y	�L�q�_�L��P�a�ĭ��l���v�����R���.���)V��|�������	z�i�j��lp���O��y����׷�����0�8�����꭭>���;���ɽ�*<e1? ��6�+t�c�K�]��s�kɽ�*<eɽ�*<eɽ�*<eY[v�_���ܑ��h"z<�'~�f7=.��ɽ�*<emD�ْ�dh89QN��hz�;3��PY���F��
�W���[�&���2�%��od�t�[.�[����V���/��!I�2�/���%�c�i�#J?�{�/z����P�V?C{u�h��@ɽ�*<e����n��r����@��և�`��$�%�ܧ�	\�j�<�U�q�Y��2�K+׷�����0yyֶ�T@�����n��..
A���ɽ�*<eNM{9q��W���P�#��6*+�'�F�W����ɽ�*<e�+�
�na���g�_Ш6�E�.8��l@�ࣨSɽ�*<e����옯��U�&4�W�{�g��"�#F��8#��U��Zv���y�1�$W.����|�TErǃ+3��|��V8��+ Z1wg�i"yPɽ�*<e8�q�ѱ�V8��+ Z��Moi��v���<���^185G��T��82�9�Sd�~�fT ��w����"vЅ\��b�]���x�\�uɽ�*<eن�\�)�e#<�޼ż�l�G��ɽ�*<e�+�
�na���g�_Zm��B��H�@�p1w�	�6�cɽ�*<e�����D��N_��^[V�Cg�����P��/���%�c�i�#J?�{�/z���"o��D�$@�՛�f��Iă�A����n��rɽ�*<e��_NN���U�ݣ��d��-QJX��~?�W#E)�dC��`E���փ<�~v3����U������h
�K=4Y[v�_�+�n�/�G��`K�f��9üI`�̸B���'�UO�����;��Y�aa24�2G7���"�#F��8����T�ҝ[��R�"`�cd �!�(I켇y��k~�G������r#��U��Z1��zfA�kC����m�@�-�F��I�|�ЮH���<���^#z�͌�?�(<��P�ay��b���4�Qp?3�w7]�'m��"�,w#��d�r"�:Dx��pɽ�*<eɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ��`���)6C�b�MPɽ�*<e-&J�� ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ곞�&`I���'d������{��Q�h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<eu;�Qݷ�2U���m)�[��/���?��a�磅"��Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<ej	�%w\������~�W%8n��Y�f�.��!I�2gː�Ï��/eJR�k�/eJR�k�/eJR�k̩�o�w
H��VJUT���	D��:�^�����%��j��\�J�����'��{
duzɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e��M�R��Lc �Ij�a�*�QW+�_�����gY��h
�K=4ɽ�*<eɽ�*<eɽ�*<eɽ�*<e����n��r�����/�\U9��8P�,[h�
�+ɽ�*<eS�;��$�Q�]�Q�Mɽ�*<eɽ�*<eɽ�*<eɽ�*<e��s��Q�V�B�f��^� |�Φ�-C��z����pɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e)�,3u�A��e6�ڡ}X}�+5��D��ݹ�Vɽ�*<e-&J�� ɽ�*<eɽ�*<eɽ�*<eɽ�*<e,4���?w��=�wYh�ǵ�\�)eE�;QC�q��i=�Z ���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<eu;�Qݷ�2U���m�|6*]�&��Jd�q/ݖ+ �0��MK�s�Zɽ�*<eɽ�*<eɽ�*<eɽ�*<ej	�%w\�����TZm��I�1�o%���G�c�тb��x���ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�VJUT���	D��:�^�����%9��z-����hԚԾ3��Q���d�O��]���/XY�-=��b��8B`}���}ͦO��/ĘsR�B�z�`u�tj&��1�����+���G:fGv�{�
;�N�s$w�h�'�h
�K=4ɽ�*<eҝ[��R��GtՑn�sW��lU%'�09k� �Nd"�O��S*��j��ΗCf�|�H蘗���?�	Qo��Q�]�Q�Mɽ�*<e�����H�*��h�A�B�R$ \�^p�!Pɽ�*<e��@�� ���q|����7#ub�^ {�Eɽ�*<e�VJUT���?�(<���JLs����٣O��Z"�#F��8�o���J|\���ֻ'��\yJ�	<�i�~��)G5�td'�b�]�������n��rɽ�*<eB��gJ��A���4�Qp?�G��q���˃�6��RbS/��~�ڭWH���.a_�A]͛Y6���K�am@��m�����x�\�uɽ�*<eن�\�)�e#<�޼����Xv�kɽ�*<e�
v�ƒm���X��cQ�]�Q�Mɽ�*<eɽ�*<eɽ�*<eҝ[��R�-��fΡ��k��4t�pԖ�����Mhɽ�*<eO��'��P�n�/ͻ�:||hy�6"pUw����^���F洰L���xr��<I}�k��b0Su���e�/���%��#��w����.�NH�h
�K=4ɽ�*<eɽ�*<e����n��r�K,V[d�@c��l2!A���K<����-�"�Y�n���[�U�~/VQPXp�P�Q�]�Q�Mɽ�*<eɽ�*<ex�\�uɽ�*<e�m=����9(�p7���������Y܄�^�7�8��إ�O�^ {�Eɽ�*<eɽ�*<eɽ�*<eY[v�_�+�n�/�G�߷G�ey2�����j���X����5�l��@�x��z>I��_jk�#��ɽ�*<eɽ�*<eɽ�*<eҝ[��R��2R&�N5݄p��P2��*�?���Y��̸B����/D��wgB��$�J�����d<��5�2-ɽ�*<eɽ�*<eNM{9q��"Rݗ]T��G5�td'�e#<�޼��+��%�ٰ���˫��5�l��@�S���B����<���^8x��*<��ɽ�*<eɽ�*<eҝ[��R���#)ϫ��K�am@��uZ1����k�I9^�ï�Lz�����K�P ��謋:��5���ڵE
\�<����(.��W��٣O��Z\�kܥ��q�/���%���7�1��kC����:���0r�=@�ࣨSɽ�*<e����n��rf3���W�����h��j��G��q���..+`��$����sb����o=$W.����|���t���M
����ɽ�*<ex�\�uɽ�*<e�m=����9l�����!7��b��M&X��~?�W#��}��N?�{�/z�:�Y�e��Q�]�Q�Mɽ�*<eY[v�_�+�n�/�G�߷G�eyc�XO�_ag�̸B���'�UO���2���K,JP�>��"�#F��8����T�ɽ�*<eҝ[��R�"`�cd �!�(I��%p>J�\������^ٰ���˫�,��T"��T�����)��~��!˃�6��Rb��33��0ɽ�*<e���������Ħ�
V8��+ ZZ�'[P�u�ɽ�*<e�/���%��8[����9(ύ��Bɽ�*<eɽ�*<eɽ�*<e����n��r�G�x9��FE�&I��}Kg��@հɽ�*<e�Y��2�K+��Qݓ˟s4�)�_π ����������'�e����Ǆ���'@�}%:�=~<���%�6��4Wj̼��(yaf��ٿ�5�l��@��a���z����.�NH�h
�K=4ɽ�*<eɽ�*<eҝ[��R���6ǝsW��lU%��~-y7ɽ�*<euJJ��pq�VcҦ>�VQPXp�P�Q�]�Q�Mɽ�*<eɽ�*<e�����H�*��h�A+c�����E��4�ɽ�*<eu5����������g�}�^ {�Eɽ�*<eɽ�*<e�VJUT���?�(<���JLs����k��b0,�o��v�/���%�P���T~��zo�_jk�#��ɽ�*<eɽ�*<e����n��rɽ�*<e�����Ez�V��]W�"�#F��8#��U��Zh��j/�\
�i��m�O�����d<��5�2-ɽ�*<e,4���?wɽ�*<e8�q�ѱ�V8��+ Zk��b0˃�6��Rb9k/�i���P���Tw�7�
�2����<���^8x��*<��ɽ�*<e����n��rɽ�*<eD$敃���q�J���
�ꈍHg�8�3�F�K2f]}v���^B%96˻�ף����
P���T�b�<���z�`u�tj&��1��[��ղ�f�!��QE����~��!W:�=����ɽ�*<eɽ�*<eҝ[��R��GtՑn�sW��lU%'�09k� �Nd"�O���l�FD�V��jU�.�LMǊ��..
A���ɽ�*<eɽ�*<e�����H�*��h�A�B�R$ \�^p�!Pɽ�*<e��w�&��^Sx=��/�:�W�Ӡ��\U�>:�ɽ�*<e�VJUT���?�(<���JLs����٣O��Z"�#F��8�o���J|���{�}f$W.����|O\�;���m�B���m���������n��rɽ�*<eB��gJ��A���4�Qp?�G��q���˃�6��Rbsw�@�u!��F{N.J?�{�/z���^��P����T�ɽ�*<ex�\�uɽ�*<eن�\�)�e#<�޼����Xv�kɽ�*<e�
v�ƒm���X��cQ�]�Q�Mɽ�*<eɽ�*<eɽ�*<eҝ[��R�-��fΡ��k��4t�pԖ�����Mhɽ�*<eO��'��P�n�/ͻ�:||hy�6"pUw����^���F洰L���xr��<I}�k��b0Su���e�/���%�P���T7���F�h+�0�ɽ�*<eɽ�*<e����n��r�K,V[d�@c��l2!A���K<����-�"�Y�n��}���麲����h���h��ɽ�*<eɽ�*<ex�\�uɽ�*<e�m=����9(�p7���������Y܄�^�7{"� L�+|�0���Ѓ��&ZReX�ɽ�*<eɽ�*<eY[v�_�+�n�/�G�߷G�ey2�����j���X����5�l��@��SwC˖�A���g�@P,͔�W�7�ɽ�*<eɽ�*<eҝ[��R��2R&�N5݄p��P2��*�?���Y��̸B����/D��wg�����y*Ȍ���\�m�B���m�����ɽ�*<eNM{9q��"Rݗ]T��G5�td'�e#<�޼��+��%�ٰ���˫��5�l��@��SwC˖�A��W���U�v��<Ϭɽ�*<eɽ�*<eҝ[��R���#)ϫ��K�am@��uZ1����k�I9^�ï�Lz�����K�P ��謋:��5���ڵE
\�<��вt���o�٣O��Z\�kܥ��q�/���%�Iή�%`��kC����:���0r�=@�ࣨSɽ�*<e����n��rf3���W�����h��j��G��q���..+`��$����sb�����x�$W.����|���t���M
����ɽ�*<ex�\�uɽ�*<e�m=����9l�����!7��b��M&X��~?�W#
j���?�{�/z�:�Y�e��Q�]�Q�Mɽ�*<eY[v�_�+�n�/�G�߷G�eyc�XO�_ag�̸B���'�UO���}%^Y[�\VJP�>��"�#F��8����T�ɽ�*<eҝ[��R�"`�cd �!�(I��%p>J�\������^ٰ���˫�,��T"�˺-H嵰. ��~��!˃�6��Rb��33��0ɽ�*<e���������Ħ�
V8��+ ZZ�'[P�u�ɽ�*<e�/���%��8[����9(ύ��Bɽ�*<eɽ�*<eɽ�*<e����n��r�G�x9��FE�&I��}Kg��@հɽ�*<e�Y��2�K+��Qݓ˟s4�)�_π ����������'�e����Ǆ���'@�}%:�=~<���%�6��4Wj̼��(yaf��ٿ�5�l��@�h�/�H���.�NH�h
�K=4ɽ�*<eɽ�*<eҝ[��R���6ǝsW��lU%��~-y7ɽ�*<euJJ��p�:�pb�VQPXp�P�Q�]�Q�Mɽ�*<eɽ�*<e�����H�*��h�A+c�����E��4�ɽ�*<eu5�����Ғ ���ƙ�^ {�Eɽ�*<eɽ�*<e�VJUT���?�(<���JLs����k��b0,�o��v�/���%�P���T�=pl?4��_jk�#��ɽ�*<eɽ�*<e����n��rɽ�*<e�����Ez�V��]W�"�#F��8#��U��Zh��j/�\
~s>B`LjP�����d<��5�2-ɽ�*<e,4���?wɽ�*<e8�q�ѱ�V8��+ Zk��b0˃�6��Rb9k/�i���P���TtWu�h����<���^8x��*<��ɽ�*<e����n��rɽ�*<eD$敃���q�J���
�ꈍHg�8�3�F�K2f]}v���^B%96˻�ף����
P���T=qM���v��z�`u�tj&��1��[��ղ�fǇz��X3�JP�>��Av�'�Bɽ�*<eɽ�*<eҝ[��R��GtՑn�sW��lU%'�09k� �Nd"�O��yh�S
cP��ry�k���~��!�AE
!�ɽ�*<eɽ�*<e�����H�*��h�A�B�R$ \�^p�!Pɽ�*<e��{Y\iqS��c�P�,�)7�1��y�����ɽ�*<e�VJUT���?�(<���JLs����٣O��Z"�#F��8�o���J|n�>�B"�kC�����&u̿1�̸B�����y���C�����n��rɽ�*<eB��gJ��A���4�Qp?�G��q���˃�6��Rbsw�@�u!�7��ɇ�F�$W.����||P����J�yϦM�|.Q�]�Q�Mx�\�uɽ�*<eن�\�)�e#<�޼����Xv�kɽ�*<e�
v�ƒm���X��cQ�]�Q�Mɽ�*<eɽ�*<eɽ�*<eҝ[��R�-��fΡ��k��4t�pԖ�����Mhɽ�*<eO��'��P�n�/ͻ�:||hy�6"pUw����^���F洰L���xr��<I}�k��b0Su���e�/���%�P���T[�tC�h+�0�ɽ�*<eɽ�*<e����n��r�K,V[d�@c��l2!A���K<����-�"�Y�n��}�����Э����h��ɽ�*<eɽ�*<ex�\�uɽ�*<e�m=����9(�p7���������Y܄�^�7���I�0���Ѓ��&ZReX�ɽ�*<eɽ�*<eY[v�_�+�n�/�G�߷G�ey2�����j���X����5�l��@���|������g�@P,͔�W�7�ɽ�*<eɽ�*<eҝ[��R��2R&�N5݄p��P2��*�?���Y��̸B����/D��wg����G���Ȍ���\�m�B���m�����ɽ�*<eNM{9q��"Rݗ]T��G5�td'�e#<�޼��+��%�ٰ���˫��5�l��@���|�����W���U�v��<Ϭɽ�*<eɽ�*<eҝ[��R���#)ϫ��K�am@��uZ1����k�I9^�ï�Lz�����K�P ��謋:��5���ڵE
\�<���E�HU�٣O��Z\�kܥ��q�/���%�|2w�e�Q��kC����:���0r�=@�ࣨSɽ�*<e����n��rf3���W�����h��j��G��q���..+`��$����sbRIꐦO�j$W.����|���t���M
����ɽ�*<ex�\�uɽ�*<e�m=����9l�����!7��b��M&X��~?�W#��	�d�?�{�/z�:�Y�e��Q�]�Q�Mɽ�*<eY[v�_�+�n�/�G�߷G�eyc�XO�_ag�̸B���'�UO��������=�JP�>��"�#F��8����T�ɽ�*<eҝ[��R�"`�cd �!�(I��%p>J�\������^ٰ���˫�yh�S
cP�^��,Fwp��~��!˃�6��Rb��33��0ɽ�*<e���������Ħ�
V8��+ ZZ�'[P�u�ɽ�*<e�/���%��8[����9(ύ��Bɽ�*<eɽ�*<eɽ�*<e����n��r�G�x9��FE�&I��}Kg��@հɽ�*<e�Y��2�K+��Qݓ˟s4�)�_π ����������'�e����Ǆ���'@�}%:�=~<���%�6��4Wj̼��(yaf��ٿ�5�l��@ɥ_S��`lH���.�NH�h
�K=4ɽ�*<eɽ�*<eҝ[��R���6ǝsW��lU%��~-y7ɽ�*<euJJ��pHW�I�ľ�VQPXp�P�Q�]�Q�Mɽ�*<eɽ�*<e�����H�*��h�A+c�����E��4�ɽ�*<eu5�����ҵ��^�'�^ {�Eɽ�*<eɽ�*<e�VJUT���?�(<���JLs����k��b0,�o��v�/���%�P���T�.�Ae�+��_jk�#��ɽ�*<eɽ�*<e����n��rɽ�*<e�����Ez�V��]W�"�#F��8#��U��Zh��j/�\
��O0�|�����d<��5�2-ɽ�*<e,4���?wɽ�*<e8�q�ѱ�V8��+ Zk��b0˃�6��Rb9k/�i���P���T�L$�z�g����<���^8x��*<��ɽ�*<e����n��rɽ�*<eD$敃���q�J���
�ꈍHg�8�3�F�K2f]}v���^B%96˻�ף����
P���T������z�`u�tj&��1��[��ղ�f�ڇ��C�JP�>��Av�'�Bɽ�*<eɽ�*<eҝ[��R��GtՑn�sW��lU%'�09k� �Nd"�O��yh�S
cP�Ɖ�D��0L��~��!�AE
!�ɽ�*<eɽ�*<e�����H�*��h�A�B�R$ \�^p�!Pɽ�*<e��{Y\iq��;�T�,�)7�1��y�����ɽ�*<e�VJUT���?�(<���JLs����٣O��Z"�#F��8�o���J|;K�Raz�kC�����&u̿1�̸B�����y���C�����n��rɽ�*<eB��gJ��A���4�Qp?�G��q���˃�6��Rbsw�@�u!�t���̌$W.����||P����J�yϦM�|.Q�]�Q�Mx�\�uɽ�*<eن�\�)�e#<�޼����Xv�kɽ�*<e�
v�ƒm���X��cQ�]�Q�Mɽ�*<eɽ�*<eɽ�*<eҝ[��R�-��fΡ��k��4t�pԖ�����Mhɽ�*<eO��'��P�n�/ͻ�:||hy�6"pUw����^���F洰L���xr��<I}�k��b0Su���e�/���%�P���T�������h+�0�ɽ�*<eɽ�*<e����n��r�K,V[d�@c��l2!A���K<����-�"�Y�n��}�������b6�H�h��ɽ�*<eɽ�*<ex�\�uɽ�*<e�m=����9(�p7���������Y܄�^�7��4�0���Ѓ��&ZReX�ɽ�*<eɽ�*<eY[v�_�+�n�/�G�߷G�ey2�����j���X����5�l��@����QkK���g�@P,͔�W�7�ɽ�*<eɽ�*<eҝ[��R��2R&�N5݄p��P2��*�?���Y��̸B����/D��wg�ߕ�)���Ȍ���\�m�B���m�����ɽ�*<eNM{9q��"Rݗ]T��G5�td'�e#<�޼��+��%�ٰ���˫��5�l��@����QkK��W���U�v��<Ϭɽ�*<eɽ�*<eҝ[��R���#)ϫ��K�am@��uZ1����k�I9^�ï�Lz�����K�P ��謋:��5���ڵE
\�<���B��*����٣O��Z\�kܥ��q�/���%󬖸3����kC����:���0r�=@�ࣨSɽ�*<e����n��rf3���W�����h��j��G��q���..+`��$����sb�ϝO�}�$W.����|���t���M
����ɽ�*<ex�\�uɽ�*<e�m=����9l�����!7��b��M&X��~?�W#|m9T�g�R?�{�/z�:�Y�e��Q�]�Q�Mɽ�*<eY[v�_�+�n�/�G�߷G�eyc�XO�_ag�̸B���'�UO���������JP�>��"�#F��8����T�ɽ�*<eҝ[��R�"`�cd �!�(I��%p>J�\������^ٰ���˫�yh�S
cP�q>��Z�.���~��!˃�6��Rb��33��0ɽ�*<e���������Ħ�
V8��+ ZZ�'[P�u�ɽ�*<e�/���%��8[����9(ύ��Bɽ�*<eɽ�*<eɽ�*<e����n��r�G�x9��FE�&I��}Kg��@հɽ�*<e�Y��2�K+��Qݓ˟s4�)�_π ����������'�e����Ǆ���'@�}%:�=~<���%�6��4Wj̼��(yaf��ٿ�5�l��@�e0�5� ����.�NH�h
�K=4ɽ�*<eɽ�*<eҝ[��R���6ǝsW��lU%��~-y7ɽ�*<euJJ��p�D����vHVQPXp�P�Q�]�Q�Mɽ�*<eɽ�*<e�����H�*��h�A+c�����E��4�ɽ�*<eu5�����҉��ܠ�Xѡ^ {�Eɽ�*<eɽ�*<e�VJUT���?�(<���JLs����k��b0,�o��v�/���%�P���T��[�����_jk�#��ɽ�*<eɽ�*<e����n��rɽ�*<e�����Ez�V��]W�"�#F��8#��U��Zh��j/�\
�d;+$�.�����d<��5�2-ɽ�*<e,4���?wɽ�*<e8�q�ѱ�V8��+ Zk��b0˃�6��Rb9k/�i���P���T��!T �����<���^8x��*<��ɽ�*<e����n��rɽ�*<eD$敃���q�J���
�ꈍHg�8�3�F�K2f]}v���^B%96˻�ף����
P���T�Ryk�vT{�z�`u�tj&��1��[��ղ�fǕpᓖC�JP�>��Av�'�Bɽ�*<eɽ�*<eҝ[��R��GtՑn�sW��lU%'�09k� �Nd"�O��yh�S
cP�����N�B��~��!�AE
!�ɽ�*<eɽ�*<e�����H�*��h�A�B�R$ \�^p�!Pɽ�*<e��{Y\iqd�������,�)7�1��y�����ɽ�*<e�VJUT���?�(<���JLs����٣O��Z"�#F��8�o���J|��f�|L�kC�����&u̿1�̸B�����y���C�����n��rɽ�*<eB��gJ��A���4�Qp?�G��q���˃�6��Rbsw�@�u!�(�2Y�ǫ$W.����||P����J�yϦM�|.Q�]�Q�Mx�\�uɽ�*<eن�\�)�e#<�޼����Xv�kɽ�*<e�
v�ƒm���X��cQ�]�Q�Mɽ�*<eɽ�*<eɽ�*<eҝ[��R�-��fΡ��k��4t�pԖ�����Mhɽ�*<eO��'��P�n�/ͻ�:||hy�6"pUw����^���F洰L���xr��<I}�k��b0Su���e�/���%�P���TWWнm��h+�0�ɽ�*<eɽ�*<e����n��r�K,V[d�@c��l2!A���K<����-�"�Y�n��}��������m��h��ɽ�*<eɽ�*<ex�\�uɽ�*<e�m=����9(�p7���������Y܄�^�7|���%
�0���Ѓ��&ZReX�ɽ�*<eɽ�*<eY[v�_�+�n�/�G�߷G�ey2�����j���X����5�l��@�B�uwo���g�@P,͔�W�7�ɽ�*<eɽ�*<eҝ[��R��2R&�N5݄p��P2��*�?���Y��̸B����/D��wg�т�Ȍ���\�m�B���m�����ɽ�*<eNM{9q��"Rݗ]T��G5�td'�e#<�޼��+��%�ٰ���˫��5�l��@�B�uwo��W���U�v��<Ϭɽ�*<eɽ�*<eҝ[��R���#)ϫ��K�am@��uZ1����k�I9^�ï�Lz�����K�P ��謋:��5���ڵE
\�<�����at�٣O��Z\�kܥ��q�/���%��/�ӄi�4�kC����:���0r�=@�ࣨSɽ�*<e����n��rf3���W�����h��j��G��q���..+`��$����sb�
T����$W.����|���t���M
����ɽ�*<ex�\�uɽ�*<e�m=����9l�����!7��b��M&X��~?�W#e���I?�{�/z�:�Y�e��Q�]�Q�Mɽ�*<eY[v�_�+�n�/�G�߷G�eyc�XO�_ag�̸B���'�UO���H���5�JP�>��"�#F��8����T�ɽ�*<eҝ[��R�"`�cd �!�(I��%p>J�\������^ٰ���˫�yh�S
cP��
��S�V��~��!˃�6��Rb��33��0ɽ�*<e���������Ħ�
V8��+ ZZ�'[P�u�ɽ�*<e�/���%��8[����9(ύ��Bɽ�*<eɽ�*<eɽ�*<e����n��r�G�x9��FE�&I��}Kg��@հɽ�*<e�Y��2�K+��Qݓ˟s4�)�_π ����������'�e����Ǆ���'@�}%:�=~<���%�6��4Wj̼��(yaf��ٿ�5�l��@�oC�K$������.�NH�h
�K=4ɽ�*<eɽ�*<eҝ[��R���6ǝsW��lU%��~-y7ɽ�*<euJJ��p�5g���VQPXp�P�Q�]�Q�Mɽ�*<eɽ�*<e�����H�*��h�A+c�����E��4�ɽ�*<eu5������#����
1͡^ {�Eɽ�*<eɽ�*<e�VJUT���?�(<���JLs����k��b0,�o��v�/���%�P���T�/T2s�*?�_jk�#��ɽ�*<eɽ�*<e����n��rɽ�*<e�����Ez�V��]W�"�#F��8#��U��Zh��j/�\
�)mh�%������d<��5�2-ɽ�*<e,4���?wɽ�*<e8�q�ѱ�V8��+ Zk��b0˃�6��Rb9k/�i���P���T%�n�iS&)���<���^8x��*<��ɽ�*<e����n��rɽ�*<eD$敃���q�J���
�ꈍHg�8�3�F�K2f]}v���^B%96˻�ף����
P���T���XN]��z�`u�tj&��1��[��ղ�f��\�m0a�JP�>��Av�'�Bɽ�*<eɽ�*<eҝ[��R��GtՑn�sW��lU%'�09k� �Nd"�O��yh�S
cP�r)1�ڹ���~��!�AE
!�ɽ�*<eɽ�*<e�����H�*��h�A�B�R$ \�^p�!Pɽ�*<e��{Y\iq*��ř%(�,�)7�1��y�����ɽ�*<e�VJUT���?�(<���JLs����٣O��Z"�#F��8�o���J|��?��B��kC�����&u̿1�̸B�����y���C�����n��rɽ�*<eB��gJ��A���4�Qp?�G��q���˃�6��Rbsw�@�u!��s7�}��$W.����||P����J�yϦM�|.Q�]�Q�Mx�\�uɽ�*<eن�\�)�e#<�޼����Xv�kɽ�*<e�
v�ƒm���X��cQ�]�Q�Mɽ�*<eɽ�*<eɽ�*<eҝ[��R�-��fΡ��k��4t�pԖ�����Mhɽ�*<eO��'��P�n�/ͻ�:||hy�6"pUw����^���F洰L���xr��<I}�k��b0Su���e�/���%�P���T8f���g�h+�0�ɽ�*<eɽ�*<e����n��r�K,V[d�@c��l2!A���K<����-�"�Y�n���g�ʿ�Ϲ��$i8��h��ɽ�*<eɽ�*<ex�\�uɽ�*<e�m=����9(�p7���������Y܄�^�7�U��_��0���Ѓ��&ZReX�ɽ�*<eɽ�*<eY[v�_�+�n�/�G�߷G�ey2�����j���X����5�l��@ɜ�(ϰ�Y����g�@P,͔�W�7�ɽ�*<eɽ�*<eҝ[��R��2R&�N5݄p��P2��*�?���Y��̸B����/D��wg>��@��8�Ȍ���\�m�B���m�����ɽ�*<eNM{9q��"Rݗ]T��G5�td'�e#<�޼��+��%�ٰ���˫��5�l��@ɜ�(ϰ�Y���W���U�v��<Ϭɽ�*<eɽ�*<eҝ[��R���#)ϫ��K�am@��uZ1����k�I9^�ï�Lz�����K�P ��謋:��5���ڵE
\�<���8oRW�$X�٣O��Z\�kܥ��q�/���%��x�#αh�kC����:���0r�=@�ࣨSɽ�*<e����n��rf3���W�����h��j��G��q���..+`��$����sbdf!п�$W.����|���t���M
����ɽ�*<ex�\�uɽ�*<e�m=����9l�����!7��b��M&X��~?�W#m��3+� �?�{�/z�:�Y�e��Q�]�Q�Mɽ�*<eY[v�_�+�n�/�G�߷G�eyc�XO�_ag�̸B���'�UO��� �D�O�h>JP�>��"�#F��8����T�ɽ�*<eҝ[��R�"`�cd �!�(I��%p>J�\������^ٰ���˫�yh�S
cP�C�6�vm���~��!˃�6��Rb��33��0ɽ�*<e���������Ħ�
V8��+ ZZ�'[P�u�ɽ�*<e�/���%��8[����9(ύ��Bɽ�*<eɽ�*<eɽ�*<e����n��r�G�x9��FE�&I��}Kg��@հɽ�*<e�Y��2�K+��Qݓ˟s4�)�_π ����������'�e����Ǆ���'@�}%:�=~<���%�6��4Wj̼��(yaf��ٿ�5�l��@�"}O���:����.�NH�h
�K=4ɽ�*<eɽ�*<eҝ[��R���6ǝsW��lU%��~-y7ɽ�*<euJJ��p���9?�YAVQPXp�P�Q�]�Q�Mɽ�*<eɽ�*<e�����H�*��h�A+c�����E��4�ɽ�*<eu5������ŃQZ1���^ {�Eɽ�*<eɽ�*<e�VJUT���?�(<���JLs����k��b0,�o��v�/���%�P���T�n[�l��s�_jk�#��ɽ�*<eɽ�*<e����n��rɽ�*<e�����Ez�V��]W�"�#F��8#��U��Zh��j/�\
2V���r������d<��5�2-ɽ�*<e,4���?wɽ�*<e8�q�ѱ�V8��+ Zk��b0˃�6��Rb9k/�i���P���T�s*���|���<���^8x��*<��ɽ�*<e����n��rɽ�*<eD$敃���q�J���
�ꈍHg�8�3�F�K2f]}v���^B%96˻�ף����
P���T =sw���z�`u�tj&��1��[��ղ�f���;��Y��#ڴ-P�h+�0�ɽ�*<eɽ�*<eҝ[��R��GtՑn�sW��lU%'�09k� �Nd"�O���+�
�na���g�_���K���$�h��ɽ�*<eɽ�*<e�����H�*��h�A�B�R$ \�^p�!Pɽ�*<e1��zfA�kC������ޔ��	3�&ZReX�ɽ�*<e�VJUT���?�(<���JLs����٣O��Z"�#F��8�o���J|�c�i�#J?�{�/z�w荦xy�cV8��+ Z�h
�K=4����n��rɽ�*<eB��gJ��A���4�Qp?�G��q���˃�6��Rbsw�@�u!�T��82�9�Sd�~�fT��9��I��5�2-ɽ�*<ex�\�uɽ�*<eن�\�)�e#<�޼����Xv�kɽ�*<e�
v�ƒm���X��cQ�]�Q�Mɽ�*<eɽ�*<eɽ�*<eҝ[��R�-��fΡ��k��4t�pԖ�����Mhɽ�*<eO��'��P�n�/ͻ�:||hy�6"pUw����^���F洰L���xr��<I}�k��b0Su���e�/���%�P���T�T�_�O�h+�0�ɽ�*<eɽ�*<e����n��r�K,V[d�@c��l2!A���K<����-�"�Y�n���g�ʿ�Ϲ�����h���h��ɽ�*<eɽ�*<ex�\�uɽ�*<e�m=����9(�p7���������Y܄�^�7��e����0���Ѓ��&ZReX�ɽ�*<eɽ�*<eY[v�_�+�n�/�G�߷G�ey2�����j���X����5�l��@�W-���zӽ��g�@P,͔�W�7�ɽ�*<eɽ�*<eҝ[��R��2R&�N5݄p��P2��*�?���Y��̸B����/D��wgQC^��oȌ���\�m�B���m�����ɽ�*<eNM{9q��"Rݗ]T��G5�td'�e#<�޼��+��%�ٰ���˫��5�l��@�W-���zӡ�W���U�v��<Ϭɽ�*<eɽ�*<eҝ[��R���#)ϫ��K�am@��uZ1���ƀVh��)��&�I��J�ѹw���[�<,]�ͻlU�� <�ZBg��jx���J���9��ɽ�*<ea�|xd����F�`�� �P1s��^!�]qɽ�*<e�jI�1�;�l-�^�� �xU�ީ�Lɽ�*<e�1q6�\
E")��ҜY;������ɽ�*<e���m#P��P��E��c�"�YZR 6�q��ɽ�*<e��S�NW�ʵ��bX�ZE^�X,6�ɽ�*<e�Д��ʝh^ӽ6Ԏm����kL	��D2�/���%��eG��Z-�]�x����g$�@ɽ�*<e8�Cc��S���Sy1�CFG�؍N�}�*MO��As��ARFd����F��#��V�l�u?�u�ɽ�*<eo"�fxK�Do?��ʌl�{����/�ӸP�[$�M�$
�$h��HfTc${[�}��
ɽ�*<e��U�ۄ��g��W���P�.a7)�ɽ�*<e�/���%�q�>%��I�l�d�t������n�0�ɽ�*<e�0Q\��DUK{r���Dj8��aڦ��ɽ�*<e�+ �0���t�Ϛ.yc&�d���^�&���5ɽ�*<e�%�G��Ŏ�&��Lc�k{�ɽ�*<e7�3]N|���p��c������� 
��(*�.�N��z�Ww���n&���鋟�v2�V��O�և�vd�Nm����r�p��3f��ɽ�*<eɽ�*<e�8����\���ֻ'�[\r�R�b���ְ��;���ɽ�*<eɽ�*<e��+�J^�Q��	�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eҝ[��R�-��fΡ��k��4t�pԖ�����Mhɽ�*<e�Y��2�K+��Qݓ˟s4�)�_π ����������'�e����Ǆ�������`둺��r�H9���G�x��W��ѥ����ɽ�*<eh��j/�\
4Wj̼��ău�Y�'ɽ�*<eɽ�*<e�VJUT����~�n�e2�h	�D�1jҮ�	�y{I�7�q]�iʳ1����h�u�B��$�J�AE
!�ɽ�*<eɽ�*<eɽ�*<eY[v�_�+�n�/�G���q���G�x��W�GZ�V�sɽ�*<eh��j/�\
}��&�rS�h
�K=4ɽ�*<eɽ�*<e�VJUT���?�(<���JLs����{Z�?����B9Hl�+s��B�"����5�l��@�x��z>I��_jk�#��ɽ�*<eɽ�*<eɽ�*<eNM{9q���ҋ\�d��6��V^�i�� N���؊��SV8��+ Zu5������!`h FH�
�̸B�����y���C�ɽ�*<eɽ�*<e�����w[i����Ç̸B���6�l�{H���R����<���^v�^7���8��إ�O�"vЅ\��b�]���ɽ�*<eɽ�*<ex�\�uɽ�*<eن�\�)�e#<�޼�.}�0/+�Su���e�/���%�\���ֻ'�[\r�R�VJ4��F���̌L�+$��9�^8�7,4���?wp�L�u*���9�k���{Z�?����}��&�rSɽ�*<e�����+���G:fGv��Y����#2��V��2�ia�s�aɽ�*<eNM{9q����Ԫ�N��iAfyl�o���ه����Jd�q/�@�j/�j��ڭWH��3�A�f<��T�;��i�.�!/O�|�*������n��rɽ�*<e�����ER�4�l�!`h FH�
�̸B���p������>�j��Ehf�+3yH&���z<�=��L�PlC�V8��+ Z�iE����n+�n�/�G�����d<��pR0N��>��7���"vЅ\��a�k|jZ�����������XPs�P2�0x����j��T�����<���^#z�͌�?�(<��P�ay��b���4�Qp?��'S�5��I>/�4	(yaf��ٿ��eRۼ����h+�0�ɽ�*<eɽ�*<eɽ�*<e}��Q�ڤ(�s:<�\��	3�Zq��2��z�..+`��"�Y�n��Z���^S��~-y7�h
�K=4ɽ�*<eɽ�*<e����n��rɽ�*<e��_NN����'S�5��u F�y��X�����eR���Z���_jk�#��ɽ�*<eɽ�*<eɽ�*<eҝ[��R��2R&�N5݄p��P2���P低ܱ"GZ�V�sɽ�*<e:��J8x���0���Ѓ��&ZReX�ɽ�*<eɽ�*<e�VJUT���?�(<���JLs����-6gɼBVzc�XO�_ag�̸B����,7�-� ����ȁĠ����d<��5�2-ɽ�*<eɽ�*<eNM{9q��"Rݗ]T��G5�td'�e#<�޼�l<��b���"vЅ\�J3�W�`>+�ݱX���+��%�yϦM�|.Q�]�Q�Mɽ�*<e,4���?wɽ�*<e�e	�5S�B���@%��,;Ԟ0��� �ɽ�*<e��@�� ���q|���afP�W���)��e�LUW:�=����ɽ�*<e&�������w=���`�M⨍ˀ��P~O�g�q]�iʳ1�Y�3�9��F�t�e�W���ߺ�i�TF�ۣ��X�Y6�M
����x�\�uɽ�*<e�m=����9��,;ԞE��4�ɽ�*<e��@�� ���q|���afP�W���)��e�LUw�	�6�cɽ�*<e����옿��P���#�l	��i�.�!/�B�"����&�JG��b�j��Ehf�+3yH&�t,�M"�Ž��g�@P,͔�W�7�Y[v�_�+�n�/�G�ƚ����'S�5��L�PlC�V8��+ ZS*��j��ΗCf�|��$EB<b eE���A�"�#F��8����T�ҝ[��R�"`�cd �!�(I�r�++����_�`/I�W6���<���^���8Yg&ڭWH��3�A�f<㋞�TUn�ñ�*�jCe�V8��+ Z�7F'�]hɽ�*<eD$敃���pR0N��>��7������P�ɽ�*<e����������XPs�P2�0x���h�@��j��{��^4�VJUT���L6�>������� +�+o��[}[��z��I-�C8�RF(Lb����(O%��;!��1�"�-�nP�[%���Q�)y�7cϢA�:��^ے���Xv�kɽ�*<eǋ'H)�@w����a���h
�K=4ɽ�*<eɽ�*<eɽ�*<eY[v�_����r�<,�����K�����]ɽ�*<e�Y��2�K+��Qݓ˟s4�)�_π ����������'�e����Ǆ�΁�K�o��c�{��%B{$A͙t�r���d��-QJ@�j/�j��ڭWH��3�A�f<��T�;��.����T�3@�ࣨS����n��r!ՠ��s����")٣O��Z��K�`ɽ�*<e����������XPs�P2�0x���o���ه���_jk�#���VJUT���?�(<��$Ǟ�2ߊ$�l�	��p�n �u�HY49�iv (�&�JG��b�j��Ehf�+3yH&���z<�=�ŏ�T��qQ�]�Q�MY[v�_�ɽ�*<e�#f̨�~��C��.���!�(I켡ֺ�e���F�t�e�W���ߺ�[�egX��Ȍ���\�m�B���*c�n��&ɽ�*<eB��gJ��A���4�Qp?�G��q���˃�6��Rb9k/�i���\���ֻ'�[\r�R�VJ4��F�����?Պl�K�am@�Z<�}U�'�ɽ�*<eP�ay��b���4�Qp?�G��q���..+`���/���%�\���ֻ'�[\r�R�VJ4��F�����r7�7}w�	�6�c,4���?w�NX�Jj�*���� )�d��\�kܥ��qɽ�*<e|�bj̜��f;��@�!W:�=����ɽ�*<eɽ�*<e�VJUT���?�(<��Vy�t�AR����Z���jME���:ɽ�*<e_'��)��_�,�\����v믜�LQ�]�Q�Mɽ�*<eɽ�*<eҝ[��R�W���P�#��6*+�'�Na(�;�49�iv (	�?�o�.�u^jP��:���Bo��h
�K=4ɽ�*<eɽ�*<eY[v�_�ɽ�*<e�#f̨�~�����J�J=��џ����	���B������
��:O�|�*��ɽ�*<eɽ�*<ex�\�uɽ�*<e�����Ez�V��]W�8�� �a�ٰ���˫��.f�nn�%ס���"�#F��8����T�ɽ�*<eɽ�*<e�����"`�cd �!�(I��%p>J�\��D�!# ٰ���˫�PI߬H��k����"V��A|m����T�ɽ�*<eɽ�*<eNM{9q��+�n�/�G˃�6��Rb�%p>J�\2����8�(yaf��ٿ�PI߬H��k�����x�����h
�K=4ɽ�*<eɽ�*<eNM{9q����X��6���`K�f^t
�`��q]�iʳ1�����	���B����Vh�jcf��Iă�Aɽ�*<eɽ�*<ex�\�uɽ�*<e��_NN��y�pn�-A�!I�2�/���%�1�"�-�ߒy�7�	�y�����ɽ�*<eɽ�*<e,4���?wɽ�*<e�JLs����[C�KZW(��K�`ɽ�*<e|�bj̜��F��y�o����7`Q�]�Q�Mɽ�*<e�VJUT���?�(<��$Ǟ�2ߊ$�l�	��p5�ε�����̸B�����͇�s6u^jP��:-̕�ո��m�B���m�����ɽ�*<eY[v�_�ɽ�*<e����o���S�B���@%!Od" [�R���<���^[�7�т����=a�^4��X�yAe�K�am@��m�����ɽ�*<e����n��rɽ�*<e�e	�5S�B���@%q�5��d��-QJw�;L�::���=a�^����y�f��9�^8�7ɽ�*<eɽ�*<e����n��r�K,V[d�"eUb^�l,�g�ǚ����P�ɽ�*<e|�bj̜��u�?[)����AE
!�ɽ�*<eɽ�*<e�VJUT���?�(<��H�*��h�A+c�����d� ��Y��ɽ�*<e_'��)��_�,�\��q�5�=�Blɽ�*<eɽ�*<eɽ�*<eҝ[��R���Ԫ�N��%/vZr���铫h���X����PI߬H��k������2�?��,͔�W�7�ɽ�*<eɽ�*<eNM{9q��+�n�/�G�ƚ������+�����d<�- �Ƈ���1�"�-U����U�G5�td'�b�]���ɽ�*<e,4���?wɽ�*<eg*D����Vm�B���Hc�ōTC���L�������of�.f�nn�]��k�hFN�"vЅ\��b�]���ɽ�*<eɽ�*<e�������#)ϫ��K�am@�Hc�ōTC�r���l&�ɽ�*<e�.f�nn��^[���ԭAv�'�Bɽ�*<eɽ�*<eɽ�*<e����영\�\R˧�sW��lU%���{K�/�Nd"�O���PI߬H��k����7�4*E(IQ�h
�K=4ɽ�*<eɽ�*<eNM{9q��+�n�/�G���q��`���o4(m������������	���B��� �[�n ���&ZReX�ɽ�*<eɽ�*<ex�\�uɽ�*<e:��8*$7���w��@����Jd�q/�w�;L�::���=a�^�A|��J�"���ɽ�*<eɽ�*<e����n��rɽ�*<e�5ŀ�@$������0*����V8��+ Z_'��)��_�,�\��xξ>�fyϦM�|.Q�]�Q�Mɽ�*<eҝ[��R�"Rݗ]T��G5�td'�e#<�޼��+�����V8��+ Z	�?�o�.�u^jP��:���(��myϦM�|.Q�]�Q�Mɽ�*<eY[v�_�ɽ�*<eن�\�)�e#<�޼�m�%���j&��1��	�?�o�.�u^jP��:&�Ջ��`
ău�Y�'ɽ�*<eɽ�*<eY[v�_����֗� q���$�*	����e�����-�w�;L�::���=a�^$��HP���h��ɽ�*<eɽ�*<e����n��rɽ�*<e�Ef�]�雈'���Y��# N��ɽ�*<e|�bj̜���`�j�Y�iw�	�6�cɽ�*<eɽ�*<e�VJUT���?�(<����P���w��(�{/U Qz�[��%�w/�.f�nn��f%*��e���K�`�h
�K=4ɽ�*<eɽ�*<e������2R&�N5݄p��P2���|C�/7&�!�(I��[��@�hk���B���l}ڞ9mx>�̸B�����y���C�ɽ�*<ex�\�uɽ�*<eB��gJ��A���4�Qp?�et�ؿ˃�6��Rb9k/�i���1�"�-9�H{L�����<���^��y���C�ɽ�*<e,4���?wɽ�*<eP�ay��b���4�Qp?�G�J,L�'Su���e�/���%�1�"�-�C�\�BPh+�0�ɽ�*<eɽ�*<e,4���?w�p\�Ì�:�C��?�^9[?y�4��}_��ɽ�*<e�.f�nn�	E�-�"u�ᦲc�ɽ�*<eɽ�*<eɽ�*<e������`���{B�3��G-}~��.�ɽ�*<e�PI߬H��k����KMFV��Q�]�Q�Mɽ�*<eɽ�*<eNM{9q��+�n�/�G�߷G�ey�a�V���>�B�"���	�?�o�.�u^jP��:����OD������ɽ�*<eɽ�*<eY[v�_�ɽ�*<e��������A���"�#F��8#��U��Z|�bj̜��ꗡ��E�������d<��5�2-ɽ�*<e�VJUT���?�(<��w[i����Ç̸B���mq�WvMEG2Ϭ%���#��U��Z_'��)��_�,�\���<sEvT�5�2-ɽ�*<eɽ�*<eҝ[��R��m�v�����<���^mq�WvMEG�$V���ɽ�*<e_'��)��_�,�\��q��̓�J�Q�]�Q�Mɽ�*<eɽ�*<eҝ[��R���s+�K���Ş��i?�lP���j�<�U�q	�?�o�.�u^jP��:&U9�Ex�M
����ɽ�*<eɽ�*<eY[v�_�ɽ�*<e�m=����9{ �ckJN��b��M&w�;L�::���=a�^t&*���	��\U�>:�ɽ�*<eɽ�*<e����n��rɽ�*<e�� Qx����0z2W��,�o��v�/���%�1�"�-o��W��_jk�#��ɽ�*<eɽ�*<e,4���?wɽ�*<e
�'63���� ~�u�zH�8��m�B�����so�[+�k����M��KV�pV8��+ Z�h
�K=4ɽ�*<eNM{9q��+�n�/�G�����d<��pR0N8��[8"[n�K�am@�*�l4h�_���B������7��w�V8��+ Z�h
�K=4ɽ�*<ex�\�uɽ�*<eD$敃���pR0NE��l�_�k��:��*ȟ����	���B������ƾ�@�ࣨSɽ�*<eɽ�*<ex�\�u�����`�
U�d	�4k"`� D..+`���/���%�1�"�-0O�P�P�..
A���ɽ�*<eɽ�*<e,4���?wɽ�*<e��K��@�W��vw�������ɽ�*<e�.f�nn�����@E��^ {�Eɽ�*<eɽ�*<eɽ�*<e����옵��������|�f�S�������G�c�т_'��)��_�,�\���� !!�ڭ�oqE�ɽ�*<eɽ�*<eҝ[��R��ҋ\�d��6��V^���c�V�G5�td'�b'��o���=a�^�6s�H����!�(I���33��0ɽ�*<e����n��rɽ�*<e8�q�ѱ�V8��+ Z�h�f����"vЅ\��a�k|jZ�|�bj̜���_P���a�˃�6��Rb��33��0ɽ�*<e�VJUT���?�(<������Ħ�
V8��+ Z�t����#\�kܥ��qɽ�*<e|�bj̜���)[���/fW:�=����ɽ�*<eɽ�*<e�VJUT���?�(<���O��3w���Z����)�`?i�ɽ�*<e_'��)��_�,�\��|I���u<�Q�]�Q�Mɽ�*<eɽ�*<eҝ[��R�W���P�#��6*+�'Й�vB�49�iv (	�?�o�.�u^jP��:'m8����h
�K=4ɽ�*<eɽ�*<eY[v�_�ɽ�*<e�#f̨�~��Fg��J�J=��џ����	���B�����qje�.0O�|�*��ɽ�*<eɽ�*<ex�\�uɽ�*<e�����Ez�V��]W���pC��v_ٰ���˫��.f�nn��/�}�|�*"�#F��8����T�ɽ�*<eɽ�*<e�����"`�cd �!�(I��%p>J�\�w�����ٰ���˫�PI߬H��k�����-4���z�����T�ɽ�*<eɽ�*<eNM{9q��+�n�/�G˃�6��Rb�%p>J�\��Wlq2"(yaf��ٿ�PI߬H��k�������N�Q�h
�K=4ɽ�*<eɽ�*<eNM{9q��gfA�q)���`K�f�e��	Q�q]�iʳ1�����	���B���ێ�L�9�f��Iă�Aɽ�*<eɽ�*<ex�\�uɽ�*<e��_NN����0��_>��!I�2�/���%�1�"�-:���n�y�����ɽ�*<eɽ�*<e,4���?wɽ�*<e�JLs����g׫��4��K�`ɽ�*<e|�bj̜�����j�� �o����7`Q�]�Q�Mɽ�*<e�VJUT���?�(<��$Ǟ�2ߊ$�l�	��p[,]!u�K;�̸B�����͇�s6u^jP��:��\(]uA�m�B���m�����ɽ�*<eY[v�_�ɽ�*<e����o���S�B���@%��'R1����<���^[�7�т����=a�^�X$�/Sn��K�am@��m�����ɽ�*<e����n��rɽ�*<e�e	�5S�B���@%똆�G�Su���ew�;L�::���=a�^(����>�h+�0�ɽ�*<eɽ�*<e����n��r�����`��"�b��jC[C�KZW(iiͱH�Rɽ�*<e|�bj̜���z_'3��ᦲc�ɽ�*<eɽ�*<e�VJUT���?�(<��H�*��h�A+c�������U>:�=�ɽ�*<e_'��)��_�,�\��#�� ���bQ�]�Q�Mɽ�*<eɽ�*<eҝ[��R���Ԫ�N��%/vZr��o��b����B�"����PI߬H��k����R��{�F��D������ɽ�*<eɽ�*<eNM{9q��+�n�/�G�ƚ��ɔ�ppJv^"�#F��8�o���J|1�"�-�U���Q�����d<��5�2-ɽ�*<e,4���?wɽ�*<eg*D����Vm�B���Hc�ōTC�|�g�� #��U��Z�.f�nn�za�^2�0}<��m��5�2-ɽ�*<eɽ�*<e�������#)ϫ��K�am@�Hc�ōTCvt8�@�Jɽ�*<e�.f�nn�za�^2�0=TS�4���Q�]�Q�Mɽ�*<eɽ�*<e�����ŵ_Dl��sW��lU%~rW蜠�k�j�<�U�q�PI߬H��k����ܦ���I��M
����ɽ�*<eɽ�*<eNM{9q��+�n�/�G���q��Z`,#�V��b��M&�����	���B�����U�=�4�\U�>:�ɽ�*<eɽ�*<ex�\�uɽ�*<e:��8*$7���I�Kw�,�o��vw�;L�::���=a�^�'�~��_jk�#��ɽ�*<eɽ�*<e����n��rɽ�*<e�5ŀ�@$�����O�3��qwm�B���hR����jD�_�,�\����"�[�V8��+ Z�h
�K=4ɽ�*<eҝ[��R�"Rݗ]T��G5�td'�e#<�޼�]��ޥ�K�am@����o��Du^jP��:C��'06�V8��+ ZL�q�e���ɽ�*<eY[v�_�ɽ�*<eن�\�)�m�H�w���9a�н�r�����׀t���8ο�K���D!�}9h����?���ג$OJ�7�/��|:��^ے���Xv�kɽ�*<eǋ'H)�@w����a���h
�K=4ɽ�*<eɽ�*<eɽ�*<eNM{9q���4����k���A�X:胮."1Do�ɽ�*<e�,��T"���`χ�a$����^�M�"�ds��R��6G�2���-l	*vQ��/�%×�˴qZ5�mq�WvMEG0��� �ɽ�*<e�F`��� ^�����h+�0�ɽ�*<eɽ�*<eɽ�*<e�������R�z����Z���l>j�m�ɽ�*<e�F`��� ^#����X�..
A���ɽ�*<eɽ�*<eɽ�*<e�����H�*��h�A+c�����E��4�ɽ�*<e�F`��� ^ ���н��y�����ɽ�*<eɽ�*<eɽ�*<e����옿��P���w��(��K�`ɽ�*<e=�i>�N�.�����UF�"���ɽ�*<eɽ�*<e�VJUT���?�(<��
�'63���� ~�u�L�PlC�V8��+ Z�PI߬H������ȁĠ����d<��5�2-ɽ�*<eɽ�*<eҝ[��R�"`�cd �!�(I��%p>J�\��W���#��U��Z�PI߬H������ȁ�˃�6��Rb��33��0ɽ�*<eɽ�*<eҝ[��R���#)ϫ��K�am@�ʮ,��7���f�}Kɽ�*<e�.f�nn�%ס���Av�'�Bɽ�*<eɽ�*<e�VJUT���ԇT^'ҵ�ۅN�����V�h�jz�i� P�ɽ�*<e�.f�nn�%ס����ᦲc�ɽ�*<eɽ�*<e�VJUT���?�(<���K��@��Y����~�|2��G�c�т�.f�nn�%ס�����K�`�h
�K=4ɽ�*<e�VJUT���?�(<��
�'63���� ~�uKlR41u49�iv (�PI߬H��k�����h=�ɗbQ�]�Q�Mɽ�*<eɽ�*<eҝ[��R����������Py�y��>��m�B���hR����jD�_�,�\��8�� �a�yϦM�|.Q�]�Q�Mɽ�*<e�����w[i����Ç̸B���i&?:�w|Gb��f	>ٰ���˫�_'��)��_�,�\��}<��m���Cה��ɽ�*<eɽ�*<e���������Ħ�
V8��+ Z+�+o��[}[��z��I-�C8�RF(Lb����(O%��;!�ٓH'b6]b=��K�XU��41�{���	����W/�6���Xv�kɽ�*<eǋ'H)�@w����a���h
�K=4ɽ�*<eɽ�*<eɽ�*<eNM{9q���4����k���A�X:胮."1Do�ɽ�*<e�,��T"���`χ�a$����^�M�"�ds��R��6G�2���-l	*vQ��/�%×�˴qZ5�mq�WvMEG0��� �ɽ�*<e�F`��� ^ .=2�����.�NH�h
�K=4ɽ�*<eɽ�*<e�������R�z����Z���l>j�m�ɽ�*<e�F`��� ^ .=2����~-y7�h
�K=4ɽ�*<eɽ�*<e�����H�*��h�A+c�����E��4�ɽ�*<e�F`��� ^ .=2��ŏ�T��qQ�]�Q�Mɽ�*<eɽ�*<e����옿��P���w��(��K�`ɽ�*<e=�i>�N���0yB�̴[���MĞ��ڭ�oqE�ɽ�*<e�VJUT���?�(<��
�'63���� ~�u�L�PlC�V8��+ Z�PI߬H���/�ʸ�}Ȍ���\�m�B���m�����ɽ�*<eҝ[��R�"`�cd �!�(I��%p>J�\��W���#��U��Z�PI߬H���/�ʸ�}�+��%�yϦM�|.Q�]�Q�Mɽ�*<eҝ[��R���#)ϫ��K�am@�ʮ,��7���f�}Kɽ�*<e�.f�nn�za�^2�0Av�'�Bɽ�*<eɽ�*<e�VJUT���ԇT^'ҵ�ۅN�����V�h�jz�i� P�ɽ�*<e�.f�nn�za�^2�0�ᦲc�ɽ�*<eɽ�*<e�VJUT���?�(<���K��@��Y����~�|2��G�c�т�.f�nn�za�^2�0��K�`�h
�K=4ɽ�*<e�VJUT���?�(<��
�'63���� ~�uKlR41u49�iv (�PI߬H��k����:�V�s

�Q�]�Q�Mɽ�*<eɽ�*<eҝ[��R����������Py�y��>��m�B���hR����jD�_�,�\��	/wx�ۻ�yϦM�|.Q�]�Q�Mɽ�*<e�����w[i����Ç̸B���i&?:�w|Gb��f	>ٰ���˫�_'��)��_�,�\���F�x�N��Cה��ɽ�*<eɽ�*<e���������Ħ�
V8��+ Z+�+o��[}[��z��I-�C8�RF(Lb����(O%��;!�ٓH'b6]b=��K�XU��41�{���	���b�<�����Xv�kɽ�*<eǋ'H)�@w����a���h
�K=4ɽ�*<eɽ�*<eɽ�*<eNM{9q���4����k���A�X:胮."1Do�ɽ�*<e�,��T"���`χ�a$����^�M�"�ds��R��6G�2���-l	*vQ��/�%×�˴qZ5�mq�WvMEG0��� �ɽ�*<e�F`��� ^
a���aF.���.�NH�h
�K=4ɽ�*<eɽ�*<e�������R�z����Z���l>j�m�ɽ�*<e�F`��� ^
a���aF.��~-y7�h
�K=4ɽ�*<eɽ�*<e�����H�*��h�A+c�����E��4�ɽ�*<e�F`��� ^
a���aF.ŏ�T��qQ�]�Q�Mɽ�*<eɽ�*<e����옿��P���w��(��K�`ɽ�*<e=�i>�N� PزK`Q[���MĞ��ڭ�oqE�ɽ�*<e�VJUT���?�(<��
�'63���� ~�u�L�PlC�V8��+ Z�PI߬H���S�B���kȌ���\�m�B���m�����ɽ�*<eҝ[��R�"`�cd �!�(I��%p>J�\��W���#��U��Z�PI߬H���S�B���k�+��%�yϦM�|.Q�]�Q�Mɽ�*<eҝ[��R���#)ϫ��K�am@�ʮ,��7���f�}Kɽ�*<e�.f�nn�]��k�hFNAv�'�Bɽ�*<eɽ�*<e�VJUT���ԇT^'ҵ�ۅN�����V�h�jz�i� P�ɽ�*<e�.f�nn�]��k�hFN�ᦲc�ɽ�*<eɽ�*<e�VJUT���?�(<���K��@��Y����~�|2��G�c�т�.f�nn�]��k�hFN��K�`�h
�K=4ɽ�*<e�VJUT���?�(<��
�'63���� ~�uKlR41u49�iv (�PI߬H��k�����h)�]�Q�]�Q�Mɽ�*<eɽ�*<eҝ[��R����������Py�y��>��m�B���hR����jD�_�,�\����_@��%yϦM�|.Q�]�Q�Mɽ�*<e�����w[i����Ç̸B���i&?:�w|Gb��f	>ٰ���˫�_'��)��_�,�\�����L����Cה��ɽ�*<eɽ�*<e���������Ħ�
V8��+ Z+�+o��[}[��z��I-�C8�RF(Lb����(O%��;!�ٓH'b6]b=��K�XU��41�{���	���C���״Y���Xv�kɽ�*<eǋ'H)�@w����a���h
�K=4ɽ�*<eɽ�*<eɽ�*<eNM{9q���4����k���A�X:胮."1Do�ɽ�*<e�,��T"���`χ�a$����^�M�"�ds��R��6G�2���-l	*vQ��/�%×�˴qZ5�mq�WvMEG0��� �ɽ�*<e�F`��� ^�Y�R�i�����.�NH�h
�K=4ɽ�*<eɽ�*<e�������R�z����Z���l>j�m�ɽ�*<e�F`��� ^�Y�R�i�⾏~-y7�h
�K=4ɽ�*<eɽ�*<e�����H�*��h�A+c�����E��4�ɽ�*<e�F`��� ^�Y�R�i��ŏ�T��qQ�]�Q�Mɽ�*<eɽ�*<e����옿��P���w��(��K�`ɽ�*<e=�i>�N�|80�2A[���MĞ��ڭ�oqE�ɽ�*<e�VJUT���?�(<��
�'63���� ~�u�L�PlC�V8��+ Z�PI߬H������d�JȌ���\�m�B���m�����ɽ�*<eҝ[��R�"`�cd �!�(I��%p>J�\��W���#��U��Z�PI߬H������d�J�+��%�yϦM�|.Q�]�Q�Mɽ�*<eҝ[��R���#)ϫ��K�am@�ʮ,��7���f�}Kɽ�*<e�.f�nn��^[���ԭAv�'�Bɽ�*<eɽ�*<e�VJUT���ԇT^'ҵ�ۅN�����V�h�jz�i� P�ɽ�*<e�.f�nn��^[���ԭ�ᦲc�ɽ�*<eɽ�*<e�VJUT���?�(<���K��@��Y����~�|2��G�c�т�.f�nn��^[���ԭ��K�`�h
�K=4ɽ�*<e�VJUT���?�(<��
�'63���� ~�uKlR41u49�iv (�PI߬H��k����V�X��Q�]�Q�Mɽ�*<eɽ�*<eҝ[��R����������Py�y��>��m�B���hR����jD�_�,�\��xξ>�fyϦM�|.Q�]�Q�Mɽ�*<e�����w[i����Ç̸B���i&?:�w|Gb��f	>ٰ���˫�_'��)��_�,�\���!��/Ϫg��Cה��ɽ�*<eɽ�*<e���������Ħ�
V8��+ Z+�+o��[}[��z��I-�C8�RF(Lb����(O%��;!�ٓH'b6]b=��K�XU��41�{���	��=qM���v����Xv�kɽ�*<eǋ'H)�@w����a���h
�K=4ɽ�*<eɽ�*<eɽ�*<eNM{9q���4����k���A�X:胮."1Do�ɽ�*<e�,��T"���`χ�a$����^�M�"�ds��R��6G�2���-l	*vQ��/�%×�˴qZ5�mq�WvMEG0��� �ɽ�*<e�F`��� ^�k�Oڴf����.�NH�h
�K=4ɽ�*<eɽ�*<e�������R�z����Z���l>j�m�ɽ�*<e�F`��� ^�k�Oڴfྏ~-y7�h
�K=4ɽ�*<eɽ�*<e�����H�*��h�A+c�����E��4�ɽ�*<e�F`��� ^�k�Oڴf�ŏ�T��qQ�]�Q�Mɽ�*<eɽ�*<e����옿��P���w��(��K�`ɽ�*<e=�i>�N��utm&Y[���MĞ��ڭ�oqE�ɽ�*<e�VJUT���?�(<��
�'63���� ~�u�L�PlC�V8��+ Z�PI߬H����%hJT7Ȍ���\�m�B���m�����ɽ�*<eҝ[��R�"`�cd �!�(I��%p>J�\��W���#��U��Z�PI߬H����%hJT7�+��%�yϦM�|.Q�]�Q�Mɽ�*<eҝ[��R���#)ϫ��K�am@�ʮ,��7���f�}Kɽ�*<e�.f�nn��f%*��e�Av�'�Bɽ�*<eɽ�*<e�VJUT���ԇT^'ҵ�ۅN�����V�h�jz�i� P�ɽ�*<e�.f�nn��f%*��e��ᦲc�ɽ�*<eɽ�*<e�VJUT���?�(<���K��@��Y����~�|2��G�c�т�.f�nn��f%*��e���K�`�h
�K=4ɽ�*<e�VJUT���?�(<��
�'63���� ~�uKlR41u49�iv (�PI߬H��k������F�Q�]�Q�Mɽ�*<eɽ�*<eҝ[��R����������Py�y��>��m�B���hR����jD�_�,�\����Y����yϦM�|.Q�]�Q�Mɽ�*<e�����w[i����Ç̸B���i&?:�w|Gb��f	>ٰ���˫�_'��)��_�,�\��OaXo�����Cה��ɽ�*<eɽ�*<e���������Ħ�
V8��+ Z+�+o��[}[��z��I-�C8�RF(Lb����(O%��;!�ٓH'b6]b=��K�XU��41�{���	����a�;Th���Xv�kɽ�*<eǋ'H)�@w����a���h
�K=4ɽ�*<eɽ�*<eɽ�*<eNM{9q���4����k���A�X:胮."1Do�ɽ�*<e�,��T"���`χ�a$����^�M�"�ds��R��6G�2���-l	*vQ��/�%×�˴qZ5�mq�WvMEG0��� �ɽ�*<e�F`��� ^!M��ch���.�NH�h
�K=4ɽ�*<eɽ�*<e�������R�z����Z���l>j�m�ɽ�*<e�F`��� ^!M��ch��~-y7�h
�K=4ɽ�*<eɽ�*<e�����H�*��h�A+c�����E��4�ɽ�*<e�F`��� ^!M��chŏ�T��qQ�]�Q�Mɽ�*<eɽ�*<e����옿��P���w��(��K�`ɽ�*<e=�i>�N��_��/�d�[���MĞ��ڭ�oqE�ɽ�*<e�VJUT���?�(<��
�'63���� ~�u�L�PlC�V8��+ Z�PI߬H����IÎȌ���\�m�B���m�����ɽ�*<eҝ[��R�"`�cd �!�(I��%p>J�\��W���#��U��Z�PI߬H����IÎ�+��%�yϦM�|.Q�]�Q�Mɽ�*<eҝ[��R���#)ϫ��K�am@�ʮ,��7���f�}Kɽ�*<e�.f�nn�	E�-�"uAv�'�Bɽ�*<eɽ�*<e�VJUT���ԇT^'ҵ�ۅN�����V�h�jz�i� P�ɽ�*<e�.f�nn�	E�-�"u�ᦲc�ɽ�*<eɽ�*<e�VJUT���?�(<���K��@��Y����~�|2��G�c�т�.f�nn�	E�-�"u��K�`�h
�K=4ɽ�*<e�VJUT���?�(<��
�'63���� ~�uKlR41u49�iv (�PI߬H��k����KMFV��Q�]�Q�Mɽ�*<eɽ�*<eҝ[��R����������Py�y��>��m�B���hR����jD�_�,�\����(�4�1�yϦM�|.Q�]�Q�Mɽ�*<e�����w[i����Ç̸B���i&?:�w|Gb��f	>ٰ���˫�_'��)��_�,�\���<sEvT��Cה��ɽ�*<eɽ�*<e���������Ħ�
V8��+ Z+�+o��[}[��z��I-�C8�RF(Lb����(O%��;!�ٓH'b6]b=��K�XU��41�{���	����������Xv�kɽ�*<eǋ'H)�@w����a���h
�K=4ɽ�*<eɽ�*<eɽ�*<eNM{9q���4����k���A�X:胮."1Do�ɽ�*<e�,��T"���`χ�a$����^�M�"�ds��R��6G�2���-l	*vQ��/�%×�˴qZ5�mq�WvMEG0��� �ɽ�*<e�F`��� ^�qֺ|*����.�NH�h
�K=4ɽ�*<eɽ�*<e�������R�z����Z���l>j�m�ɽ�*<e�F`��� ^�qֺ|*Ӿ�~-y7�h
�K=4ɽ�*<eɽ�*<e�����H�*��h�A+c�����E��4�ɽ�*<e�F`��� ^�qֺ|*�ŏ�T��qQ�]�Q�Mɽ�*<eɽ�*<e����옿��P���w��(��K�`ɽ�*<e=�i>�N�lC�z�q�[���MĞ��ڭ�oqE�ɽ�*<e�VJUT���?�(<��
�'63���� ~�u�L�PlC�V8��+ Z�PI߬H��o,�)Nk�Ȍ���\�m�B���m�����ɽ�*<eҝ[��R�"`�cd �!�(I��%p>J�\��W���#��U��Z�PI߬H��o,�)Nk��+��%�yϦM�|.Q�]�Q�Mɽ�*<eҝ[��R���#)ϫ��K�am@�ʮ,��7���f�}Kɽ�*<e�.f�nn�+�2���Av�'�Bɽ�*<eɽ�*<e�VJUT���ԇT^'ҵ�ۅN�����V�h�jz�i� P�ɽ�*<e�.f�nn�+�2����ᦲc�ɽ�*<eɽ�*<e�VJUT���?�(<���K��@��Y����~�|2��G�c�т�.f�nn�+�2�����K�`�h
�K=4ɽ�*<e�VJUT���?�(<��
�'63���� ~�uKlR41u49�iv (�PI߬H��k�����<dtFnQ�]�Q�Mɽ�*<eɽ�*<eҝ[��R����������Py�y��>��m�B���hR����jD�_�,�\���q�0g�yϦM�|.Q�]�Q�Mɽ�*<e�����w[i����Ç̸B���i&?:�w|Gb��f	>ٰ���˫�_'��)��_�,�\��{x�e�6���Cה��ɽ�*<eɽ�*<e���������Ħ�
V8��+ Z+�+o��[}[��z��I-�C8�RF(Lb����(O%��;!�ٓH'b6]b=��K�XU��41�{���	��J��a����Xv�kɽ�*<eǋ'H)�@w����a���h
�K=4ɽ�*<eɽ�*<eɽ�*<eNM{9q���4����k���A�X:胮."1Do�ɽ�*<e�,��T"���`χ�a$����^�M�"�ds��R��6G�2���-l	*vQ��/�%×�˴qZ5�mq�WvMEG0��� �ɽ�*<e�F`��� ^���������.�NH�h
�K=4ɽ�*<eɽ�*<e�������R�z����Z���l>j�m�ɽ�*<e�F`��� ^�����ʾ�~-y7�h
�K=4ɽ�*<eɽ�*<e�����H�*��h�A+c�����E��4�ɽ�*<e�F`��� ^������ŏ�T��qQ�]�Q�Mɽ�*<eɽ�*<e����옿��P���w��(��K�`ɽ�*<e=�i>�N��d�����I[���MĞ��ڭ�oqE�ɽ�*<e�VJUT���?�(<��
�'63���� ~�u�L�PlC�V8��+ Z�PI߬H��n<ˋ�DMȌ���\�m�B���m�����ɽ�*<eҝ[��R�"`�cd �!�(I��%p>J�\��W���#��U��Z�PI߬H��n<ˋ�DM�+��%�yϦM�|.Q�]�Q�Mɽ�*<eҝ[��R���#)ϫ��K�am@�ʮ,��7���f�}Kɽ�*<e�.f�nn�����@E�Av�'�Bɽ�*<eɽ�*<e�VJUT���ԇT^'ҵ�ۅN�����V�h�jz�i� P�ɽ�*<e�.f�nn�����@E��ᦲc�ɽ�*<eɽ�*<e�VJUT���?�(<���K��@��Y����~�|2��G�c�т�.f�nn�����@E���K�`�h
�K=4ɽ�*<e�VJUT���?�(<��
�'63���� ~�uKlR41u49�iv (�PI߬H��k������(W �vQ�]�Q�Mɽ�*<eɽ�*<eҝ[��R����������Py�y��>��m�B���hR����jD�_�,�\���>���c�yϦM�|.Q�]�Q�Mɽ�*<e�����w[i����Ç̸B���i&?:�w|Gb��f	>ٰ���˫�_'��)��_�,�\�����3\����Cה��ɽ�*<eɽ�*<e���������Ħ�
V8��+ Z+�+o��[}[��z��I-�C8�RF(Lb����(O%��;!�ٓH'b6]b=��K�XU��41�{���	���Ryk�vT{���Xv�kɽ�*<eǋ'H)�@w����a���h
�K=4ɽ�*<eɽ�*<eɽ�*<eNM{9q���4����k���A�X:胮."1Do�ɽ�*<e�,��T"���`χ�a$����^�M�"�ds��R��6G�2���-l	*vQ��/�%×�˴qZ5�mq�WvMEG0��� �ɽ�*<e�F`��� ^�yC�~|5���.�NH�h
�K=4ɽ�*<eɽ�*<e�������R�z����Z���l>j�m�ɽ�*<e�F`��� ^�yC�~|5��~-y7�h
�K=4ɽ�*<eɽ�*<e�����H�*��h�A+c�����E��4�ɽ�*<e�F`��� ^�yC�~|5ŏ�T��qQ�]�Q�Mɽ�*<eɽ�*<e����옿��P���w��(��K�`ɽ�*<e=�i>�N�Z�I�]�4[���MĞ��ڭ�oqE�ɽ�*<e�VJUT���?�(<��
�'63���� ~�u�L�PlC�V8��+ Z�PI߬H����RzLPȌ���\�m�B���m�����ɽ�*<eҝ[��R�"`�cd �!�(I��%p>J�\��W���#��U��Z�PI߬H����RzLP�+��%�yϦM�|.Q�]�Q�Mɽ�*<eҝ[��R���#)ϫ��K�am@�ʮ,��7���f�}Kɽ�*<e�.f�nn��/�}�|�*Av�'�Bɽ�*<eɽ�*<e�VJUT���ԇT^'ҵ�ۅN�����V�h�jz�i� P�ɽ�*<e�.f�nn��/�}�|�*�ᦲc�ɽ�*<eɽ�*<e�VJUT���?�(<���K��@��Y����~�|2��G�c�т�.f�nn��/�}�|�*��K�`�h
�K=4ɽ�*<e�VJUT���?�(<��
�'63���� ~�uKlR41u49�iv (�PI߬H��k�����v����N�Q�]�Q�Mɽ�*<eɽ�*<eҝ[��R����������Py�y��>��m�B���hR����jD�_�,�\����pC��v_yϦM�|.Q�]�Q�Mɽ�*<e�����w[i����Ç̸B���i&?:�w|Gb��f	>ٰ���˫�_'��)��_�,�\���"�����Cה��ɽ�*<eɽ�*<e���������Ħ�
V8��+ Z+�+o��[}[��z��I-�C8�RF(Lb����(O%��;!�ٓH'b6]b=��K�XU��41�{���	��y��	�ϣ����Xv�kɽ�*<eǋ'H)�@w����a���h
�K=4ɽ�*<eɽ�*<eɽ�*<eNM{9q���4����k���A�X:胮."1Do�ɽ�*<e�,��T"���`χ�a$����^�M�"�ds��R��6G�2���-l	*vQ��/�%×�˴qZ5�mq�WvMEG0��� �ɽ�*<e�F`��� ^\ѯ
��?����.�NH�h
�K=4ɽ�*<eɽ�*<e�������R�z����Z���l>j�m�ɽ�*<e�F`��� ^\ѯ
��?���~-y7�h
�K=4ɽ�*<eɽ�*<e�����H�*��h�A+c�����E��4�ɽ�*<e�F`��� ^\ѯ
��?�ŏ�T��qQ�]�Q�Mɽ�*<eɽ�*<e����옿��P���w��(��K�`ɽ�*<e=�i>�N���0>)�k�[���MĞ��ڭ�oqE�ɽ�*<e�VJUT���?�(<��
�'63���� ~�u�L�PlC�V8��+ Z�PI߬H���q �y�Ȍ���\�m�B���m�����ɽ�*<eҝ[��R�"`�cd �!�(I��%p>J�\��W���#��U��Z�PI߬H���q �y��+��%�yϦM�|.Q�]�Q�Mɽ�*<eҝ[��R���#)ϫ��K�am@�ʮ,��7���f�}Kɽ�*<e�.f�nn��W6����\Av�'�Bɽ�*<eɽ�*<e�VJUT���ԇT^'ҵ�ۅN�����V�h�jz�i� P�ɽ�*<e�.f�nn��W6����\�ᦲc�ɽ�*<eɽ�*<e�VJUT���?�(<���K��@��Y����~�|2��G�c�т�.f�nn��W6����\��K�`�h
�K=4ɽ�*<e�VJUT���?�(<��
�'63���� ~�uKlR41u49�iv (�PI߬H��k����`1�JQ��SQ�]�Q�Mɽ�*<eɽ�*<eҝ[��R����������Py�y��>��m�B���hR����jD�_�,�\����D8QXz�yϦM�|.Q�]�Q�Mɽ�*<e�����w[i����Ç̸B���i&?:�w|Gb��f	>ٰ���˫�_'��)��_�,�\��t�99�`���Cה��ɽ�*<eɽ�*<e���������Ħ�
V8��+ Z+�+o��[}[��z��I-�C8�RF(Lb����(O%��;!�ٓH'b6]b=��K�XU��41�{���	�����XN]����Xv�kɽ�*<eǋ'H)�@w����a���h
�K=4ɽ�*<eɽ�*<eɽ�*<eNM{9q���4����k���A�X:胮."1Do�ɽ�*<e�,��T"���`χ�a$����^�M�"�ds��R��6G�2���-l	*vQ��/�%×�˴qZ5�mq�WvMEG0��� �ɽ�*<e�F`��� ^W�nS�?����.�NH�h
�K=4ɽ�*<eɽ�*<e�������R�z����Z���l>j�m�ɽ�*<e�F`��� ^W�nS�?���~-y7�h
�K=4ɽ�*<eɽ�*<e�����H�*��h�A+c�����E��4�ɽ�*<e�F`��� ^W�nS�?�ŏ�T��qQ�]�Q�Mɽ�*<eɽ�*<e����옿��P���w��(��K�`ɽ�*<e=�i>�N��6�$?��[���MĞ��ڭ�oqE�ɽ�*<e�VJUT���?�(<��
�'63���� ~�u�L�PlC�V8��+ Z�PI߬H��9�5P,�Ȍ���\�m�B���m�����ɽ�*<eҝ[��R�"`�cd �!�(I��%p>J�\��W���#��U��Z�PI߬H��9�5P,��+��%�yϦM�|.Q�]�Q�Mɽ�*<eҝ[��R���#)ϫ��K�am@�ʮ,��7���f�}Kɽ�*<e�.f�nn�za�^2�0<�%K\�d�Q�]�Q�Mɽ�*<e�VJUT���ԇT^'ҵ�ۅN�����V�h�jz�i� P�ɽ�*<e�.f�nn�za�^2�0��v믜�LQ�]�Q�Mɽ�*<e�VJUT���?�(<���K��@��Y����~�|2��G�c�т�.f�nn�za�^2�0�8����c��ڭ�oqE�ɽ�*<e�VJUT���?�(<��
�'63���� ~�uKlR41u49�iv (�PI߬H��k������U>:�=��h
�K=4ɽ�*<eɽ�*<eҝ[��R����������Py�y��>��m�B���hR����jD�_�,�\��U�V�]�$V8��+ Z�h
�K=4ɽ�*<e�����w[i����Ç̸B���i&?:�w|Gb��f	>ٰ���˫�_'��)��_�,�\���|�g�� U�v��<Ϭɽ�*<eɽ�*<e���������Ħ�
V8��+ Z+�+o��[}[��z��I-�C8�RF(Lb����(O%��;!�ٓH'b6]b=��K�XU��41�{���	���o���D�i���Xv�kɽ�*<eǋ'H)�@w����a���h
�K=4ɽ�*<eɽ�*<eɽ�*<eNM{9q���4����k���A�X:胮."1Do�ɽ�*<e�,��T"���`χ�a$����^�M�"�ds��R��6G�2���-l	*vQ��/�%×�˴qZ5�mq�WvMEG0��� �ɽ�*<e�F`��� ^�lx�������.�NH�h
�K=4ɽ�*<eɽ�*<e�������R�z����Z���l>j�m�ɽ�*<e�F`��� ^�lx���þ�~-y7�h
�K=4ɽ�*<eɽ�*<e�����H�*��h�A+c�����E��4�ɽ�*<e�F`��� ^�lx����ŏ�T��qQ�]�Q�Mɽ�*<eɽ�*<e����옿��P���w��(��K�`ɽ�*<e=�i>�N�Vnl�@�2�[���MĞ��ڭ�oqE�ɽ�*<e�VJUT���?�(<��
�'63���� ~�u�L�PlC�V8��+ Z�PI߬H��n!B�dYoȌ���\�m�B���m�����ɽ�*<eҝ[��R�"`�cd �!�(I��%p>J�\��W���#��U��Z�PI߬H��n!B�dYo�+��%�yϦM�|.Q�]�Q�Mɽ�*<eҝ[��R���#)ϫ��K�am@�ʮ,��7���f�}Kɽ�*<e�.f�nn�za�^2�0=TS�4���Q�]�Q�Mɽ�*<e�VJUT���ԇT^'ҵ�ۅN�����V�h�jz�i� P�ɽ�*<e�.f�nn�za�^2�0�=߂���Q�]�Q�Mɽ�*<e�VJUT���?�(<���K��@��Y����~�|2��G�c�т�.f�nn�za�^2�0�aE������ڭ�oqE�ɽ�*<e�VJUT���?�(<��
�'63���� ~�uKlR41u49�iv (�PI߬H��k�����tJe�����h
�K=4ɽ�*<eɽ�*<eҝ[��R����������Py�y��>��m�B���hR����jD�_�,�\����"�[�V8��+ Z�h
�K=4ɽ�*<e�����w[i����Ç̸B���i&?:�w|Gb��f	>ٰ���˫�_'��)��_�,�\��V�I��@�U�v��<Ϭɽ�*<eɽ�*<e���������Ħ�
V8��+ Z+�+o��[}[��z��I-�C8�RF(Lb����(O%��;!���E��!��nP�[%���Q�)y��|P�:��^ے���Xv�kɽ�*<e�
v�ƒm���X��cQ�]�Q�Mɽ�*<eɽ�*<eɽ�*<eҝ[��R�-��fΡ��k��4t�pԖ�����Mhɽ�*<eO��'��P�n�/ͻ�:||hy�6"pUw����^���F洰L���xr��<I}�٣O��Z\�kܥ��q�/���%�P���T���c�h+�0�ɽ�*<eɽ�*<e����n��rf3���W�����h��j��G��q���,�o��v"�Y�n��}����"��'L��Σ"���ɽ�*<eɽ�*<ex�\�uɽ�*<e������٣O��ZY��# N���/���%�P���T8����y�����ɽ�*<eɽ�*<e����n��rɽ�*<e:��8*$7��.m`.t�G5�td'��S#n0ŧ|j�����!`h FH�
�̸B�����y���C�ɽ�*<eY[v�_�+�n�/�G�����d<��pR0N/�Z8�{��K�am@����H�fd;��z�*�+��%�yϦM�|.Q�]�Q�Mɽ�*<eNM{9q���m�v�����<���^i&?:�w� b��ɽ�*<eu5����������g�}�ᦲc�ɽ�*<eɽ�*<e�VJUT���?�(<���K��@�W��vw!����� �ɽ�*<e,F���u_%f;��@�!W:�=����ɽ�*<eɽ�*<e,4���?w�K,V[d��*���/w)�d������P��/���%��E��!��
��)k�j..
A���ɽ�*<eɽ�*<e����n��rɽ�*<e��_NN��I���~L�=�!I�2"�Y�n���t�2M�����@�^��\U�>:�ɽ�*<eɽ�*<ex�\�uɽ�*<e�#f̨�~�����J�J=����(�ܼ�ԕu^jP��:�;������D������ɽ�*<eɽ�*<eNM{9q���ҋ\�d��6��V^���.L�G5�td'�,|	����i�~R�}ɻ�&lc�̸B�����y���C�ɽ�*<eY[v�_�+�n�/�G�����d<��pR0N�9��>֑2�K�am@������ �u^jP��:��D�!# yϦM�|.ɽ�*<eɽ�*<eNM{9q���m�v�����<���^��5��ޝt�=	E���;�V�
%��
Y\�er"�꺯z^��>��q����?���ג$OJ�7��d�cF):�k�P˥̹尮l;�DhY��F�ɽ�*<e��=!��(2��p�ɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���MO�~Iy'p�k�ɽ�*<e$����sb����o=�����bC�x���b��6�-4�)�_π۷9�V$�K�o��c�{��%B{$A͙t�r���d��-QJ�Y܄�^�7{"� L�+|.����T�3@�ࣨSɽ�*<eɽ�*<eY[v�_�J3�"�K���`K�f� �C�ZJ�J=��ѫ���h�u������y*2�����j�D������ɽ�*<eɽ�*<eNM{9q���ҋ\�d��6��V^�l�����!7��b��M&�Y܄�^�7{"� L�+|�0���Ѓ��&ZReX�ɽ�*<eɽ�*<eY[v�_�+�n�/�G�߷G�eyc�XO�_ag�̸B����I�?4ز�SwC˖�A�L�PlC�V8��+ Z�h
�K=4ɽ�*<eҝ[��R�"`�cd �!�(I��%p>J�\������^ٰ���˫�uJJ��p{3"Xf)�u���v��{�5�2-ɽ�*<eɽ�*<e���������Ħ�
V8��+ Z٣O��Z����P��/���%�P���T���ãņ..
A���ɽ�*<eɽ�*<e����n��rɽ�*<e��_NN��I���~L�=Su���e"�Y�n���t�2M�����g�}<�%K\�d�Q�]�Q�Mɽ�*<ex�\�uv�L{Ǘ%>���$�*���~PS����-����~�I���i�~R�۷��Y��ᦲc�ɽ�*<eɽ�*<eY[v�_�+�n�/�G���q��3�f�>7���������(�ܼ�ԕ��02v6cS&�*;w�	�6�cɽ�*<eɽ�*<eNM{9q����Ԫ�N��%/vZr���;��������X�����>�A�%�k�P˥-�{����"���ɽ�*<eɽ�*<e�����$Ǟ�2ߊ$�l�	��p�}ɻ�&lc�̸B����,7�-� �⧼��-�z߷7��1sG5�td'�b�]���ɽ�*<eҝ[��R�"`�cd �!�(I��%p>J�\��D�!# ٰ���˫��>�A�%�k�P˥��>?��'��K�am@���QX�T�>ɽ�*<e���������Ħ�
V8��+ Z+�+o��[}[��z��I-�C8�RF(Lb����(O%��;!���E��!��nP�[%���Q�)y��|P��K��G�,BZ�'[P�u�ɽ�*<e�/���%��8[����9(ύ��Bɽ�*<eɽ�*<eɽ�*<e����n��r�G�x9��FE�&I��}Kg��@հɽ�*<e�Y��2�K+��Qݓ˟s4�)�_π ����������'�e����Ǆ���'@�}%:�=~<���%�6���z�`u�tj&��1���5�l��@�h�/�H���.�NH�h
�K=4ɽ�*<eɽ�*<eҝ[��R��GtՑn�sW��lU%�u F�y��X���uJJ��p�:�pb�[���MĞ��ڭ�oqE�ɽ�*<eɽ�*<e�����$Ǟ�2ߊ$�l�	��p�n �u�HY49�iv (�5�l��@�h�/�Hŏ�T��qQ�]�Q�Mɽ�*<eɽ�*<eҝ[��R����������Py��؊��SV8��+ Zu5�����Ғ ���ƙ"�#F��8����T�ɽ�*<e�VJUT���?�(<��g*D����Vm�B���ʮ,��7�|M��t+c�����ofh��j/�\
~s>B`LjP˃�6��Rb��33��0ɽ�*<e,4���?wɽ�*<e�e	�5S�B���@%C�xW�a����-��Y܄�^�7wڤBRWd��ٰ#sf��Iă�Aɽ�*<eɽ�*<eY[v�_�+�n�/�G���q�������'��:��*��(�ܼ�ԕ��02v6c�p�s W:�=����ɽ�*<eɽ�*<eNM{9q��Z',`�Á��Ş��i$�EC���j�<�U�q)ԙ=Llm6�⧼��-����>��..
A���ɽ�*<eɽ�*<eҝ[��R��`���{B�3��G���Bo�ɽ�*<e��>�A�%�R��+�����@�^��\U�>:�ɽ�*<eɽ�*<e����옿��P���w��(�8����c�[��%�w/,F���u_%
a���aF.�;������D������ɽ�*<e,4���?wɽ�*<e�5ŀ�@$�����+)��S�*5V8��+ Z�k�O�O�S�B���k�}ɻ�&lc�̸B�����y���C��VJUT���?�(<��g*D����Vm�B���Hc�ōTC}<��m������of,F���u_%
a���aF.��D�!# yϦM�|.ɽ�*<e,4���?wɽ�*<e�e	�5S�B���@%9��z-����hԚԾ3��Q���d�O��]�㮇en�^^����i�~Rb=��K�X�y�]�eC�t�2M�5����w��'ѳ��w��ɽ�*<e1? ��6�+t�c�K�]��s�kɽ�*<eɽ�*<eɽ�*<eY[v�_���ܑ��h"z<�'~�f7=.��ɽ�*<e�,��T"���`χ�a$����^�M�"�ds��R��6G�2���-l	*vQ��/�%×�˴qZ5�i&?:�w������ɽ�*<eu5������i?�����)Av�'�Bɽ�*<eɽ�*<e�VJUT���n5�e֐2�h	����V�h�j��BSҧ�[��%�w/h��j/�\
��CVD�o����7`Q�]�Q�Mɽ�*<e,4���?wɽ�*<e�5ŀ�@$n���Ā�^p�!Pɽ�*<eu5������i?�����)�^ {�Eɽ�*<eɽ�*<e�VJUT���?�(<���JLs����٣O��Z"�#F��8�o���J|P���T�z0� xG5�td'�b�]���ɽ�*<e����n��rɽ�*<eB��gJ��A���4�Qp?�G��q���˃�6��Rbd�*���j}����\���}u@�K�am@��m�����ɽ�*<ex�\�uɽ�*<eن�\�)�e#<�޼�}!�Lڜ�j�<�U�q�5�l��@���|�����~-y7�h
�K=4ɽ�*<eɽ�*<eҝ[��R��`���{B�3��G旿�]��(yaf��ٿ��>�A�%ӿ�F��+ �Q� _9���9�^8�7ɽ�*<eɽ�*<e�����Vy�t�AR����Z���jME���:ɽ�*<e�k�O�O����d�J$�EC��f��Iă�Aɽ�*<e�VJUT���?�(<���K��@�W��vw#
%��+�ɽ�*<e,F���u_%�Y�R�i�����Bo��h
�K=4ɽ�*<e,4���?wɽ�*<e�� Qx���I���~L�=,�o��v"�Y�n���t�2M�� ���ƙ�8����c��ڭ�oqE�ɽ�*<ex�\�uɽ�*<e������)�d��"�#F��8�o���J|�E��!�|80�2A+)��S�*5V8��+ Z�h
�K=4����n��rɽ�*<eB��gJ��A���4�Qp?I���~L�=˃�6��Rbd�*���j�t�2M�� ���ƙ}<��m���Cה��ɽ�*<ex�\�uɽ�*<eن�\�)�m�H�w���9a�н�r�����׀t���8ο�K����Xq��wˆ㯪�@��]�ͻlU��	��	�����02v6c=qM���v����Xv�kɽ�*<e�
v�ƒm���X��cQ�]�Q�Mɽ�*<eɽ�*<eɽ�*<eҝ[��R�-��fΡ��k��4t�pԖ�����Mhɽ�*<eO��'��P�n�/ͻ�:||hy�6"pUw����^���F洰L���xr��<I}�٣O��Z\�kܥ��q�/���%�P���T�jwQy��h+�0�ɽ�*<eɽ�*<e����n��rf3���W�����h��j��G��q���,�o��v"�Y�n��}���麪Öl�u�4�"���ɽ�*<eɽ�*<ex�\�uɽ�*<e������٣O��ZY��# N���/���%�P���T���i#�y�����ɽ�*<eɽ�*<e����n��rɽ�*<e:��8*$7��.m`.t�G5�td'��S#n0�B9X�N���!`h FH�
�̸B�����y���C�ɽ�*<eY[v�_�+�n�/�G�����d<��pR0N/�Z8�{��K�am@����H�fCz���U%�+��%�yϦM�|.Q�]�Q�Mɽ�*<eNM{9q���m�v�����<���^i&?:�w� b��ɽ�*<eu5�����ҵ��^�'�ᦲc�ɽ�*<eɽ�*<e�VJUT���?�(<���K��@�W��vw!����� �ɽ�*<e,F���u_%�k�Oڴf�旿�]��ău�Y�'ɽ�*<e,4���?w�K,V[d��*���/w)�d������P��/���%��E��!��utm&YjME���:�h
�K=4ɽ�*<e����n��rɽ�*<e��_NN��I���~L�=�!I�2"�Y�n���t�2M�i?�����)2�1D���ɽ�*<eɽ�*<ex�\�uɽ�*<e�#f̨�~�����J�J=����(�ܼ�ԕ��02v6c�H1dȿ��o����7`Q�]�Q�Mɽ�*<eNM{9q���ҋ\�d��6��V^���.L�G5�td'�,|	����i�~R(��z�ƣ"�#F��8����T�ɽ�*<eY[v�_�+�n�/�G�����d<��pR0N�9��>֑2�K�am@������ ���02v6c�H1dȿ�˃�6��Rb�8dY�֚
ɽ�*<eNM{9q���m�v�����<���^��5��ޝt�=	E���;�V�
%��
Y\�er"�꺯z^��>��q����?���ג$OJ�7��d�cF):����>>�̹尮l;�DhY��F�ɽ�*<e��=!��(2��p�ɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���MO�~Iy'p�k�ɽ�*<e$����sb����o=�����bC�x���b��6�-4�)�_π۷9�V$�K�o��c�{��%B{$A͙t�r���d��-QJ�Y܄�^�7��4.����T�3@�ࣨSɽ�*<eɽ�*<eY[v�_�J3�"�K���`K�f� �C�ZJ�J=��ѫ���h�u��ߕ�)���2�����j�D������ɽ�*<eɽ�*<eNM{9q���ҋ\�d��6��V^�l�����!7��b��M&�Y܄�^�7��4�0���Ѓ��&ZReX�ɽ�*<eɽ�*<eY[v�_�+�n�/�G�߷G�eyc�XO�_ag�̸B����I�?4ز���QkK�L�PlC�V8��+ Z�h
�K=4ɽ�*<eҝ[��R�"`�cd �!�(I��%p>J�\������^ٰ���˫�uJJ��p;�}�qn2#���v��{�5�2-ɽ�*<eɽ�*<e���������Ħ�
V8��+ Z٣O��Z����P��/���%�P���T��^-���..
A���ɽ�*<eɽ�*<e����n��rɽ�*<e��_NN��I���~L�=Su���e"�Y�n���t�2M����^�'<�%K\�d�Q�]�Q�Mɽ�*<ex�\�uv�L{Ǘ%>���$�*���~PS����-����~�I���i�~R��A��,I�ᦲc�ɽ�*<eɽ�*<eY[v�_�+�n�/�G���q��3�f�>7���������(�ܼ�ԕ��02v6c�c�f�E��w�	�6�cɽ�*<eɽ�*<eNM{9q����Ԫ�N��%/vZr���;��������X�����>�A�%����>>�-�{����"���ɽ�*<eɽ�*<e�����$Ǟ�2ߊ$�l�	��p�}ɻ�&lc�̸B����,7�-� �⧼��-�u���Ω�G5�td'�b�]���ɽ�*<eҝ[��R�"`�cd �!�(I��%p>J�\��D�!# ٰ���˫��>�A�%����>>���>?��'��K�am@���QX�T�>ɽ�*<e���������Ħ�
V8��+ Z+�+o��[}[��z��I-�C8�RF(Lb����(O%��;!���E��!��nP�[%���Q�)y��|P�H�e���}Z�'[P�u�ɽ�*<e�/���%��8[����9(ύ��Bɽ�*<eɽ�*<eɽ�*<e����n��r�G�x9��FE�&I��}Kg��@հɽ�*<e�Y��2�K+��Qݓ˟s4�)�_π ����������'�e����Ǆ���'@�}%:�=~<���%�6���z�`u�tj&��1���5�l��@�e0�5� ����.�NH�h
�K=4ɽ�*<eɽ�*<eҝ[��R��GtՑn�sW��lU%�u F�y��X���uJJ��p�D����vH[���MĞ��ڭ�oqE�ɽ�*<eɽ�*<e�����$Ǟ�2ߊ$�l�	��p�n �u�HY49�iv (�5�l��@�e0�5� �ŏ�T��qQ�]�Q�Mɽ�*<eɽ�*<eҝ[��R����������Py��؊��SV8��+ Zu5�����҉��ܠ�X�"�#F��8����T�ɽ�*<e�VJUT���?�(<��g*D����Vm�B���ʮ,��7�|M��t+c�����ofh��j/�\
�d;+$�.˃�6��Rb��33��0ɽ�*<e,4���?wɽ�*<e�e	�5S�B���@%C�xW�a����-��Y܄�^�70 A��!Md��ٰ#sf��Iă�Aɽ�*<eɽ�*<eY[v�_�+�n�/�G���q�������'��:��*��(�ܼ�ԕ��02v6c�1쀺T�W:�=����ɽ�*<eɽ�*<eNM{9q��Z',`�Á��Ş��i$�EC���j�<�U�q)ԙ=Llm6�⧼��-�N����hA..
A���ɽ�*<eɽ�*<eҝ[��R��`���{B�3��G���Bo�ɽ�*<e��>�A�%|�>��~����@�^��\U�>:�ɽ�*<eɽ�*<e����옿��P���w��(�8����c�[��%�w/,F���u_%�qֺ|*��;������D������ɽ�*<e,4���?wɽ�*<e�5ŀ�@$�����+)��S�*5V8��+ Z�k�O�Oo,�)Nk��}ɻ�&lc�̸B�����y���C��VJUT���?�(<��g*D����Vm�B���Hc�ōTC}<��m������of,F���u_%�qֺ|*ә�D�!# yϦM�|.ɽ�*<e,4���?wɽ�*<e�e	�5S�B���@%9��z-����hԚԾ3��Q���d�O��]�㮇en�^^����i�~Rb=��K�X�y�]�eC�t�2M�j��z�%e7'ѳ��w��ɽ�*<e1? ��6�+t�c�K�]��s�kɽ�*<eɽ�*<eɽ�*<eY[v�_���ܑ��h"z<�'~�f7=.��ɽ�*<e�,��T"���`χ�a$����^�M�"�ds��R��6G�2���-l	*vQ��/�%×�˴qZ5�i&?:�w������ɽ�*<eu5������Je�G%LnAv�'�Bɽ�*<eɽ�*<e�VJUT���n5�e֐2�h	����V�h�j��BSҧ�[��%�w/h��j/�\
{��S�~�o����7`Q�]�Q�Mɽ�*<e,4���?wɽ�*<e�5ŀ�@$n���Ā�^p�!Pɽ�*<eu5������Je�G%Ln�^ {�Eɽ�*<eɽ�*<e�VJUT���?�(<���JLs����٣O��Z"�#F��8�o���J|P���T��I�>EA�G5�td'�b�]���ɽ�*<e����n��rɽ�*<eB��gJ��A���4�Qp?�G��q���˃�6��Rbd�*���j}����-f��`I��K�am@��m�����ɽ�*<ex�\�uɽ�*<eن�\�)�e#<�޼�}!�Lڜ�j�<�U�q�5�l��@�B�uwo��~-y7�h
�K=4ɽ�*<eɽ�*<eҝ[��R��`���{B�3��G旿�]��(yaf��ٿ��>�A�%� Բ��+�Q� _9���9�^8�7ɽ�*<eɽ�*<e�����Vy�t�AR����Z���jME���:ɽ�*<e�k�O�On<ˋ�DM$�EC��f��Iă�Aɽ�*<e�VJUT���?�(<���K��@�W��vw#
%��+�ɽ�*<e,F���u_%���������Bo��h
�K=4ɽ�*<e,4���?wɽ�*<e�� Qx���I���~L�=,�o��v"�Y�n���t�2M����ܠ�Xџ8����c��ڭ�oqE�ɽ�*<ex�\�uɽ�*<e������)�d��"�#F��8�o���J|�E��!��d�����I+)��S�*5V8��+ Z�h
�K=4����n��rɽ�*<eB��gJ��A���4�Qp?I���~L�=˃�6��Rbd�*���j�t�2M����ܠ�X�}<��m���Cה��ɽ�*<ex�\�uɽ�*<eن�\�)�m�H�w���9a�н�r�����׀t���8ο�K����Xq��wˆ㯪�@��]�ͻlU��	��	�����02v6c�Ryk�vT{���Xv�kɽ�*<e�
v�ƒm���X��cQ�]�Q�Mɽ�*<eɽ�*<eɽ�*<eҝ[��R�-��fΡ��k��4t�pԖ�����Mhɽ�*<eO��'��P�n�/ͻ�:||hy�6"pUw����^���F洰L���xr��<I}�٣O��Z\�kܥ��q�/���%�P���TrQ�t7<�h+�0�ɽ�*<eɽ�*<e����n��rf3���W�����h��j��G��q���,�o��v"�Y�n��}�������I:T��"���ɽ�*<eɽ�*<ex�\�uɽ�*<e������٣O��ZY��# N���/���%�P���Tp ��)����y�����ɽ�*<eɽ�*<e����n��rɽ�*<e:��8*$7��.m`.t�G5�td'��S#n0�sKh��dT!`h FH�
�̸B�����y���C�ɽ�*<eY[v�_�+�n�/�G�����d<��pR0N/�Z8�{��K�am@����H�f�{l��E�_�+��%�yϦM�|.Q�]�Q�Mɽ�*<eNM{9q���m�v�����<���^i&?:�w� b��ɽ�*<eu5������#����
1��ᦲc�ɽ�*<eɽ�*<e�VJUT���?�(<���K��@�W��vw!����� �ɽ�*<e,F���u_%�yC�~|5旿�]��ău�Y�'ɽ�*<e,4���?w�K,V[d��*���/w)�d������P��/���%��E��!�Z�I�]�4jME���:�h
�K=4ɽ�*<e����n��rɽ�*<e��_NN��I���~L�=�!I�2"�Y�n���t�2M�Je�G%Ln2�1D���ɽ�*<eɽ�*<ex�\�uɽ�*<e�#f̨�~�����J�J=����(�ܼ�ԕ��02v6cP��
h�o����7`Q�]�Q�Mɽ�*<eNM{9q���ҋ\�d��6��V^���.L�G5�td'�,|	����i�~RT3�'Y�U"�#F��8����T�ɽ�*<eY[v�_�+�n�/�G�����d<��pR0N�9��>֑2�K�am@������ ���02v6cP��
h˃�6��Rb�8dY�֚
ɽ�*<eNM{9q���m�v�����<���^��5��ޝt�=	E���;�V�
%��
Y\�er"�꺯z^��>��q����?���ג$OJ�7��d�cF):L2�*<*S�̹尮l;�DhY��F�ɽ�*<e��=!��(2��p�ɽ�*<eɽ�*<eɽ�*<e�VJUT���?�(<���MO�~Iy'p�k�ɽ�*<e$����sb����o=�����bC�x���b��6�-4�)�_π۷9�V$�K�o��c�{��%B{$A͙t�r���d��-QJ�Y܄�^�7�U��_�.����T�3@�ࣨSɽ�*<eɽ�*<eY[v�_�J3�"�K���`K�f� �C�ZJ�J=��ѫ���h�u�>��@��8�2�����j�D������ɽ�*<eɽ�*<eNM{9q���ҋ\�d��6��V^�l�����!7��b��M&�Y܄�^�7�U��_��0���Ѓ��&ZReX�ɽ�*<eɽ�*<eY[v�_�+�n�/�G�߷G�eyc�XO�_ag�̸B����I�?4ز��(ϰ�Y��L�PlC�V8��+ Z�h
�K=4ɽ�*<eҝ[��R�"`�cd �!�(I��%p>J�\������^ٰ���˫�uJJ��p$�GK�a���v��{�5�2-ɽ�*<eɽ�*<e���������Ħ�
V8��+ Z٣O��Z����P��/���%�P���Tv����;..
A���ɽ�*<eɽ�*<e����n��rɽ�*<e��_NN��I���~L�=Su���e"�Y�n���t�2M�#����
1�<�%K\�d�Q�]�Q�Mɽ�*<ex�\�uv�L{Ǘ%>���$�*���~PS����-����~�I���i�~R��g+��q�ᦲc�ɽ�*<eɽ�*<eY[v�_�+�n�/�G���q��3�f�>7���������(�ܼ�ԕ��02v6c#z�C-���w�	�6�cɽ�*<eɽ�*<eNM{9q����Ԫ�N��%/vZr���;��������X�����>�A�%L2�*<*S�-�{����"���ɽ�*<eɽ�*<e�����$Ǟ�2ߊ$�l�	��p�}ɻ�&lc�̸B����,7�-� �⧼��-�}�KF@�	G5�td'�b�]���ɽ�*<eҝ[��R�"`�cd �!�(I��%p>J�\��D�!# ٰ���˫��>�A�%L2�*<*S���>?��'��K�am@���QX�T�>ɽ�*<e���������Ħ�
V8��+ Z+�+o��[}[��z��I-�C8�RF(Lb����(O%��;!���E��!��nP�[%���Q�)y��|P�9�6`BHZ�'[P�u�ɽ�*<e�/���%��8[����9(ύ��Bɽ�*<eɽ�*<eɽ�*<e����n��r�G�x9��FE�&I��}Kg��@հɽ�*<e�Y��2�K+��Qݓ˟s4�)�_π ����������'�e����Ǆ���'@�}%:�=~<���%�6���z�`u�tj&��1���5�l��@�"}O���:����.�NH�h
�K=4ɽ�*<eɽ�*<eҝ[��R��GtՑn�sW��lU%�u F�y��X���uJJ��p���9?�YA[���MĞ��ڭ�oqE�ɽ�*<eɽ�*<e�����$Ǟ�2ߊ$�l�	��p�n �u�HY49�iv (�5�l��@�"}O���:�ŏ�T��qQ�]�Q�Mɽ�*<eɽ�*<eҝ[��R����������Py��؊��SV8��+ Zu5������ŃQZ1��"�#F��8����T�ɽ�*<e�VJUT���?�(<��g*D����Vm�B���ʮ,��7�|M��t+c�����ofh��j/�\
2V���r�˃�6��Rb��33��0ɽ�*<e,4���?wɽ�*<e�e	�5S�B���@%C�xW�a����-��Y܄�^�7D�Ɂ�p��d��ٰ#sf��Iă�Aɽ�*<eɽ�*<eY[v�_�+�n�/�G���q�������'��:��*��(�ܼ�ԕ��02v6c�
�m���*W:�=����ɽ�*<eɽ�*<eNM{9q��Z',`�Á��Ş��i$�EC���j�<�U�q)ԙ=Llm6`m�J�dOn=�Ԯb�..
A���ɽ�*<eɽ�*<eҝ[��R��`���{B�3��G���Bo�ɽ�*<e��>�A�%�d-0�Ų����@�^��\U�>:�ɽ�*<eɽ�*<e����옿��P���w��(�8����c�[��%�w/,F���u_%W�nS�?��;������D������ɽ�*<e,4���?wɽ�*<e�5ŀ�@$�����+)��S�*5V8��+ Z�k�O�O9�5P,��}ɻ�&lc�̸B�����y���C��VJUT���?�(<��g*D����Vm�B���Hc�ōTC}<��m������of,F���u_%W�nS�?���D�!# yϦM�|.ɽ�*<e,4���?wɽ�*<e�e	�5S�B���@%9��z-����hԚԾ3��Q���d�O��]�㮇en�^^����i�~Rb=��K�X�y�]�eC�t�2M������Y\'ѳ��w��ɽ�*<e1? ��6�+t�c�K�]��s�kɽ�*<eɽ�*<eɽ�*<eY[v�_���ܑ��h"z<�'~�f7=.��ɽ�*<e�,��T"���`χ�a$����^�M�"�ds��R��6G�2���-l	*vQ��/�%×�˴qZ5�i&?:�w������ɽ�*<eu5������Yk�!��>Av�'�Bɽ�*<eɽ�*<e�VJUT���n5�e֐2�h	����V�h�j��BSҧ�[��%�w/h��j/�\
8�'	ϛ�i�o����7`Q�]�Q�Mɽ�*<e,4���?wɽ�*<e�5ŀ�@$n���Ā�^p�!Pɽ�*<eu5������Yk�!��>�^ {�Eɽ�*<eɽ�*<e�VJUT���?�(<���JLs����٣O��Z"�#F��8�o���J|P���TӰO/��9G5�td'�b�]���ɽ�*<e����n��rɽ�*<eB��gJ��A���4�Qp?�G��q���˃�6��Rbd�*���j�g�ʿ�Ϲ-ڲ�TrM��K�am@��m�����ɽ�*<ex�\�uɽ�*<eن�\�)�e#<�޼�}!�Lڜ�j�<�U�q�5�l��@�W-���zӾ�~-y7�h
�K=4ɽ�*<eɽ�*<eҝ[��R��`���{B�3��G旿�]��(yaf��ٿ��>�A�%��J���׌Q� _9���9�^8�7ɽ�*<eɽ�*<e�����Vy�t�AR����Z���jME���:ɽ�*<e�k�O�On!B�dYo$�EC��f��Iă�Aɽ�*<e�VJUT���?�(<���K��@�W��vw#
%��+�ɽ�*<e,F���u_%�lx�������Bo��h
�K=4ɽ�*<e,4���?wɽ�*<e�� Qx���I���~L�=,�o��v"�Y�n���t�2M�ŃQZ1���8����c��ڭ�oqE�ɽ�*<ex�\�uɽ�*<e������)�d��"�#F��8�o���J|�E��!�Vnl�@�2�+)��S�*5V8��+ Z�h
�K=4����n��rɽ�*<eB��gJ��A���4�Qp?I���~L�=˃�6��Rbd�*���j�t�2M�ŃQZ1��}<��m���Cה��ɽ�*<ex�\�uɽ�*<eن�\�)�m�H�w���9a�н�r�����׀t���8ο�K����Xq��w�����?���ג$OJ�7�Gw#x9�):��^ے���Xv�kɽ�*<e1? ��6�+t�c�K�]��s�kɽ�*<eɽ�*<eɽ�*<eY[v�_���ܑ��h"z<�'~�f7=.��ɽ�*<e�Y��2�K+��Qݓ˟s4�)�_π ����������'�e����Ǆ���'@�}%:�=~<���%�6��4Wj̼��(yaf��ٿ���~�Im��3sxL5�M�k/Q�]�Q�Mɽ�*<eɽ�*<eY[v�_��;�헳쳤`K�f����<}�j�<�U�q"�Y�n��Z���^S��~-y7�h
�K=4ɽ�*<eɽ�*<ex�\�uɽ�*<e�m=����9(�p7���������/���%��ݱX��}��&�rS�h
�K=4ɽ�*<eɽ�*<e����n��rɽ�*<e:��8*$7�~D(qza�J�J=����/���%��ݱX��2�����j�D������ɽ�*<eɽ�*<e����n��rɽ�*<e�����Ez�V��]W�"�#F��8#��U��Z��eR�&_��b��{G5�td'�b�]���ɽ�*<eɽ�*<e�����w[i����Ç̸B���mq�WvMEG���v��{�����of)ԙ=Llm6����ȁ�˃�6��Rb��33��0ɽ�*<eɽ�*<eҝ[��R���#)ϫ��K�am@�ʮ,��7���f�}Kɽ�*<e��>�A�%�_�,�\��<�%K\�d�Q�]�Q�Mɽ�*<eɽ�*<e���2��3��H�=<1>�2�04�}�1�|�0cNd"�O��)ԙ=Llm6k����jME���:�h
�K=4ɽ�*<eɽ�*<eҝ[��R��`���{B�3��G��2K�c,�B�"����(�ܼ�ԕu^jP��:�;������D������ɽ�*<eɽ�*<eNM{9q���ҋ\�d��6��V^���7�4[i�!I�2�/���%��E��!�	�����ұ�y�����ɽ�*<eɽ�*<e����n��rɽ�*<e:��8*$7���7�4[i�����d<�- �Ƈ����E��!��ߡ����G5�td'�b�]���ɽ�*<e����n��rɽ�*<eB��gJ��A���4�Qp?Nf�^)��"vЅ\��a�k|jZ�,F���u_%f;��@�!˃�6��Rb��33��0ɽ�*<e,4���?wɽ�*<e�e	�5S�B���@%(��N�lWASu���e�/���%��E��!���0yB�̴>������h
�K=4ɽ�*<e����n��rpH[��V�^��)��K�+�������P�ɽ�*<e,F���u_% .=2��py<��֋M
����ɽ�*<e,4���?wɽ�*<e�Ef�]�٣O��Z�aE�����[��%�w/�k�O�O�/�ʸ�}���
��:O�|�*��ɽ�*<e�VJUT���?�(<��
�'63���� ~�u��_�l�B49�iv (�(�ܼ�ԕ��02v6cS&�*;w�	�6�cɽ�*<eɽ�*<eNM{9q����Ԫ�N��%/vZr��iC�ͫ�U��̸B����F#��8 ��02v6cS&�*;�����d<��5�2-ɽ�*<eNM{9q��"Rݗ]T��G5�td'�e#<�޼��OG����`�K�am@��`v�C����i�~R�۷��Y��"vЅ\��b�]���ɽ�*<eY[v�_�+�n�/�G˃�6��Rb�%p>J�\iy���K�Xj&��1���(�ܼ�ԕ��02v6c�p�s W:�=����ɽ�*<eɽ�*<eNM{9q�����#Φ3g���Ş��i��>-����q]�iʳ1���~�I���i�~R�Q�����ᦲc�ɽ�*<eɽ�*<eY[v�_�+�n�/�G���q��'(ܢ��B���Jd�q/�"�Y�n���t�2M�c�A�`Pꞟ8����c��ڭ�oqE�ɽ�*<ex�\�uɽ�*<e������٣O��ZR2�*�H|Yɽ�*<e�k�O�O�S�B���k�Na(�;��&ZReX�ɽ�*<e�VJUT���?�(<���JLs����٣O��Z��_@��%ٰ���˫��k�O�O�S�B���k�}ɻ�&lc�̸B�����y���C��VJUT���?�(<��g*D����Vm�B���ʮ,��7�j�F��F,�#��U��Z��>�A�%�R��+���>?��'��K�am@��m�����ɽ�*<e���������Ħ�
V8��+ Z٣O��Z�r���l&�ɽ�*<e�k�O�O����d�J����t�@�ࣨSɽ�*<e�VJUT���ԇT^'�n�F^�� g���V�h�j�8(���=ɽ�*<e��>�A�%ӿ�F��+ ��) �)x�h��ɽ�*<eɽ�*<e�����H�*��h�A�B�R$ \q��$�F
��X���)ԙ=Llm6�⧼��-��N3��ޘ'�_jk�#��ɽ�*<eɽ�*<eҝ[��R��2R&�N5݄p��P2��X*E��!��b��M&"�Y�n���t�2M�� ���ƙ2�1D���ɽ�*<eɽ�*<ex�\�uɽ�*<e�#f̨�~h��g֧�G5�td'/O�&�Na�t�2M�� ���ƙ8�� �a�yϦM�|.Q�]�Q�Mx�\�uɽ�*<e����o���S�B���@%�6>M��:�˃�6��Rb9k/�i����E��!�|80�2A"V��A|m����T�ɽ�*<e����n��rɽ�*<eD$敃���pR0Noj��Pĝ�d��-QJ"�Y�n���t�2M�i?�����)<�%K\�d�Q�]�Q�Mɽ�*<ex�\�uc������$�*�����..+`���/���%��E��!��utm&YjME���:�h
�K=4ɽ�*<e����n��rɽ�*<e��_NN��o�,
j�F:��K�`ɽ�*<e,F���u_%�k�Oڴf��;������D������ɽ�*<e,4���?wɽ�*<e�5ŀ�@$n���Ā��"�<�ɽ�*<e)ԙ=Llm6�⧼��-��R���3 �y�����ɽ�*<eɽ�*<eҝ[��R����������Py�=kpjg���m�B���>����b��⧼��-�B��@�Y��G5�td'�b�]���ɽ�*<eҝ[��R�"`�cd �!�(I��%p>J�\���Ͳ�WV8��+ Z�(�ܼ�ԕ��02v6c�H1dȿ�˃�6��Rb��33��0ɽ�*<eNM{9q���m�v�����<���^i&?:�w������o(yaf��ٿ)ԙ=Llm6�⧼��-���識Y�ch+�0�ɽ�*<eɽ�*<eҝ[��R��c���)��sW��lU%=��m:u;�j�<�U�q�(�ܼ�ԕ��02v6c�c�f�E���AE
!�ɽ�*<eɽ�*<eNM{9q��W���P�#��6*+�'h��>T�9�J�J=��х��~�I���i�~R��A��,I��K�`�h
�K=4ɽ�*<eY[v�_�+�n�/�G�ƚ�읳#>�V��Y��# N��ɽ�*<e,F���u_%!M��ch���Bo��h
�K=4ɽ�*<e,4���?wɽ�*<e�� Qx��ӳ#>�V��"�#F��8#��U��Z,F���u_%!M��ch�[�-o�m�B���m�����,4���?wɽ�*<e8�q�ѱ�V8��+ Z٣O��Z�<sEvT�����of�k�O�O��IÎ>5xW�V8��+ Z�h
�K=4�VJUT���?�(<��P�ay��b���4�Qp?�NW1(�!X\�kܥ��qɽ�*<e,F���u_%�qֺ|*�旿�]��ău�Y�'ɽ�*<e,4���?wf3���W��K����B٣O��Z~�<+���ɽ�*<e�k�O�Oo,�)Nk�$�EC��f��Iă�Aɽ�*<e�VJUT���?�(<���K��@��Y����#��+��G�c�т��>�A�%|�>��~-�{����"���ɽ�*<eɽ�*<e�����$Ǟ�2ߊ$�l�	��p�n�Y�s�S����������~�I���i�~R���Dk�x�^ {�Eɽ�*<eɽ�*<eY[v�_�+�n�/�G�߷G�eyBtw�;���!�(I�q���D�$���i�~R���Dk�x"�#F��8����T�ɽ�*<eY[v�_�+�n�/�G�����d<��pR0N�{5��~���<���^����O�t�2M�s��ĵ��&}<��m��5�2-ɽ�*<ex�\�uɽ�*<eن�\�)�e#<�޼Ÿ�z4#R
��:��*ȅ��~�I���i�~R�l���Av�'�Bɽ�*<eɽ�*<eY[v�_��ϧY4����`K�f��!�4	�٦���-�"�Y�n���t�2M����ܠ�Xі�v믜�LQ�]�Q�Mɽ�*<ex�\�uɽ�*<e�m=����9�p��
J,�o��v�/���%��E��!��d�����I3�Q���,͔�W�7�ɽ�*<e����n��rɽ�*<e�����E1Y"�7&��В�J콷ɽ�*<e��>�A�%� Բ��+����@�^��\U�>:�ɽ�*<eɽ�*<e����옿��P����_5��휽]�����V8��+ Z��>�A�%� Բ��+���'B[t;�!�(I���33��0ɽ�*<e�����w[i����Ç̸B���i&?:�w�X�k�9.�ٰ���˫�)ԙ=Llm6�⧼��-����jP����<���^��y���C�ɽ�*<eҝ[��R���#)ϫ��K�am@�ʮ,��7��x�Gᑻɽ�*<e��>�A�%s�(��|�Q� _9���9�^8�7ɽ�*<eɽ�*<e���2��3tR��m֡2�04��L\[���Nd"�O��)ԙ=Llm6�⧼��-��y"6,��..
A���ɽ�*<eɽ�*<eҝ[��R��`���{B�3��G�j���:�'�B�"����(�ܼ�ԕ��02v6cP��
h�o����7`Q�]�Q�Mɽ�*<eNM{9q���ҋ\�d��6��V^��i\�Oک�!I�2�/���%��E��!�Z�I�]�4�h=�ɗbQ�]�Q�Mɽ�*<e����n��rɽ�*<e:��8*$7��i\�Oک�����d<�- �Ƈ����E��!�Z�I�]�4+)��S�*5V8��+ Z�h
�K=4����n��rɽ�*<eB��gJ��A���4�Qp?\��}���"vЅ\��a�k|jZ�,F���u_%�yC�~|5��D�!# yϦM�|.Q�]�Q�M,4���?wɽ�*<e�e	�5S�B���@%J��x6��[Su���e�/���%��E��!���0>)�k�>������h
�K=4ɽ�*<e����n��rpH[��V��%	=���W��׶1����P�ɽ�*<e,F���u_%\ѯ
��?�py<��֋M
����ɽ�*<e,4���?wɽ�*<e�Ef�]�٣O��Z����XC[��%�w/�k�O�O�q �y����
��:O�|�*��ɽ�*<e�VJUT���?�(<��
�'63���� ~�u���}��49�iv (�(�ܼ�ԕ��02v6c#z�C-���w�	�6�cɽ�*<eɽ�*<eNM{9q����Ԫ�N��%/vZr������� �g�̸B����F#��8 ��02v6c#z�C-�� ����d<��5�2-ɽ�*<eNM{9q��"Rݗ]T��G5�td'�e#<�޼šseFxG&��K�am@��`v�C����i�~R��g+��q�"vЅ\��b�]���ɽ�*<eY[v�_�+�n�/�G˃�6��Rb�%p>J�\�6'�05���:��*��(�ܼ�ԕ��02v6c�
�m���*W:�=����ɽ�*<eɽ�*<eNM{9q��*�!�#}�Ş��i̻���
����-����~�I���i�~R�GU_np���ᦲc�ɽ�*<eɽ�*<eY[v�_�+�n�/�G���q����#��˗,�o��v"�Y�n���t�2M��� �Oट8����c��ڭ�oqE�ɽ�*<ex�\�uɽ�*<e������٣O��Z��"׀\ɽ�*<e�k�O�O9�5P,��Na(�;��&ZReX�ɽ�*<e�VJUT���?�(<���JLs����٣O��ZU�V�]�$V8��+ Z�k�O�O9�5P,��}ɻ�&lc�̸B�����y���C��VJUT���?�(<��g*D����Vm�B���ʮ,��7����� O��ٰ���˫��>�A�%�d-0�Ų��>?��'��K�am@��m�����ɽ�*<e���������Ħ�
V8��+ Z٣O��Zvt8�@�Jɽ�*<e�k�O�On!B�dYo����t�@�ࣨSɽ�*<e�VJUT���GӼ�*�O�.$�3�<����V�h�jˌ�����PNd"�O����>�A�%��J������) �)x�h��ɽ�*<eɽ�*<e�����H�*��h�A�B�R$ \##����X �B�"���)ԙ=Llm6`m�J�ddU�i��_jk�#��ɽ�*<eɽ�*<eҝ[��R��2R&�N5݄p��P2��!�� ��!I�2"�Y�n���t�2M�ŃQZ1��2�1D���ɽ�*<eɽ�*<ex�\�uɽ�*<e�#f̨�~�!�� ˠ����d<�=c$��[�t�2M�ŃQZ1��8�� �a�yϦM�|.Q�]�Q�Mx�\�uɽ�*<e����o���S�B���@%@��}(���"vЅ\�J3�W�`>+�E��!�Vnl�@�2�"V��A|mU�v��<Ϭɽ�*<e����n��rɽ�*<eD$敃���q�J���
�ꈍHg�8�3�F�K2f]}v���^B%aj�l�t�v2}&�@B1Y-�q f�&��������r=9xϞ�(��<�uO�%�t$�!P�N�Ě̆$�>qg�\XQH����c��~/^�"�dI��sZ��w4�v�Ѽ��B�.�Xz�ϥ�l<�S�v�Ѽc�oK�SK��4ȹ�5�v�Ѽݾ!-��<���K�v�Ѽ�N�Ƴ�+ �0���v�Ѽ`��(D�+ �0���v�Ѽޞ����VǛ
}���V����Jj�|Ĳ)�48lZ��_�E�+��43nb>�����Ϡ�����|;�NF��׈�`�%�����\#�@�]mp���V�B$g�Brh�!**��NF��׈�T٫��#�Z[��� ]mp���+ ���=��v���%�]mp����kB�]$l����A�%�jF���l�ʶ�"OA%�2`�i�طt�"���l�w�a0�u,.姎��a���h
�K=4ɽ�*<eɽ�*<eɽ�*<e6��/�нf���10
����3,����;��	Զ����Qݓ˟s4�)�_π ����������'�e����ǄU���B(�{hԡj���	P�T����)���KS�$����sb����o=$W.����|c� k�k��L�����`w�	�6�cx�\�uJ�fMw~�(�߷G�ey�q�ɚ G�Z[��� ��7�1��kC����^��N2�{�&�����ڧ�ᦲc�����n��rɽ�*<e�m=����9қ�u;`J�d��-QJmD�ْ�Ad ݰm�H/��+�ͼ�f���9TI���.�NH�����?�(<����t5��;��̲�E6�#
%��+��@�v;�z���v����c5U�2#��))��h
�K=4ɽ�*<e'a���ˑ�#+�m�� �^[V�Cg�)�rj��+c�m<>�m�^�v2}&�[}ͣ��T��f�f��Iă�Aɽ�*<eNM{9q���`���{�"M��
�/"���S�|����/�]�찴�}0�@Z���ŗ<�䴗�.�h+�0�ɽ�*<ex�\�u+�n�/�G��`K�f���6��o��МB\'��ɏu��7)��S�c�Y�=��}*.�ɽ�*<e,4���?wɽ�*<e&9��? ��9q:Xx3���^������eX�3%7|P���ޤ�]�찴�}0�@Z���ŗb��i���sX!�	�u>�o��P���� /"|�"�~���G>y�[]��ɺ��L]=�����6����_Ĳ�w�P � ��jY�q���36.^�d��%YC^2����ߐuX�q�0&�r�2����-���D�ߐuX�q�Dy秤_����RG�:O�ߐuX�q�$�s~e	Ӽ�j�<�U�q}���5�lv�G�0���j&��1��}���5�l��D�.��J ��u���ߐuX�q�RDk�,$�	��-���D�~�g2H� �c��Q�S������k�d��Ję��Jߌ���%�THM�%�G��ن������H��̞d��JęXq�!x�^����-��%�G���%`���yʏd��-QJ�%�G���\
|J:�Gk]91Ŗ��8����g�����6��o�����"�dJŭ쀏D�b+f���H�����+�J^�Q��	�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��,r�/�MeN�q�Xߣ�k �y����L�>��2��`χ�a$����^�M�"�ds��R��6G�2���-l	*v��I�,��؅��U>ɺ���V���/�#
%��+��Y��2�K+ҫ�0�7Ӑ����3e�X�Bh�W�0���Ѓ��&ZReX�NM{9q���\~C����jN�̓��)�rj��+cX��~?�W#-KB�i�Sd�~�fT�[V�`��zǙ�7��h��Y[v�_�W���P�#��6*+�'��^Ii6Q�v���%����{�}f$W.����|c� k�k��L�����`W:�=��������n��rɽ�*<e���$�*�0.�#�d�!I�2dE�0(|�:B�2ƍ�zCd;��z�*8�����}�\U�>:��VJUT���y�=R)��}�����\$��I8�����P�\_*X�#~v'�w�֬����K��NJ��� ..
A���ɽ�*<e����옝�K��@��@��U��&�}�m<>�m�^�v2}&�PZ�n.{{�xq�`��Av�'�Bɽ�*<eNM{9q��!�T9�k����S��N�y��^C���w�]�찴�}0�@Z���ŗh^�g%B�#zI�-�k�L�q�e���x�\�u+�n�/�G�YN�F�N�ꈍHg�8�3�F�K2f]}v���^B%aj�l�t�v2}&�@B1Y-�q f�&��������r=9xϞ�(��<�uO�%�t$�!P�N�Ě̆$�>qg�\XQH����c��~/^�"�dI��sZ��w4�v�Ѽ��B�.�Xz�ϥ�l<�S�v�Ѽc�oK�SK��4ȹ�5�v�Ѽݾ!-��<���K�v�Ѽ�N�Ƴ�+ �0���v�Ѽ`��(D�+ �0���v�Ѽޞ����VǛ
}���V����Jj�|Ĳ)�48lZ��_�E�+��43nb>�����Ϡ�����|;�NF��׈�`�%�����\#�@�]mp���V�B$g�Brh�!**��NF��׈�T٫��#�Z[��� ]mp���+ ���=��v���%�]mp����kB�]$l����A�%�jF���l�ʶ���u�[��B{#Jĭ�B
pfo����H�R�g��1-P��V]��%�ɽ�*<eɽ�*<eɽ�*<e,4���?w�+�ږ�F�X��X�+�)�ڙ�c �_`�ͨ�O��'��P�n�/ͻ�:||hy�6"pUw����^���F洰�-_ɪ�
a��1D��7�#J.�5�!I�2�,��T"�˺-H嵰. ���W�X��<R|=-}��&�rS�h
�K=4�&�;!��l�����k��-inh����P�[��ղ�f�}%^Y[�\V�����3e�X�Bh�Wd��ٰ#sf��Iă�Aҝ[��R�H�*��h�A�5B�	��U��&�}X��~?�W#
j���?�{�/z�p�^(]e��C�]�Nf��h+�0�Y[v�_��H��g澁��Ş��i8�����}�"C�g�����6��o����k���ҿy��))��h
�K=4����n��rj9PՂ�{�#f̨�~����������-��ɏu��7)��S�Y-�m`n��f�f��Iă�A,4���?wɽ�*<e��_NN��\$��I8�\�kܥ��q\_*X�#~v'�w�֬���3��U��
<�䴗�.�h+�0�ɽ�*<e�������]/߷�W6�v����zI�-�k��m<>�m�^�v2}&�PZ�n.{{LZ�"""����}*.�ɽ�*<eNM{9q���ܡ�,�'�%=��CTZ� g�+�����ʠ��6�L�d�[s�	�4�ڟ�}�}�(�L+'�w�֬��_�1��Ø��8B`}�FW,P��/b&�'�}�����֩�*��x`E%�N��|d$o���7�3]N|�F�j�!f��=oX�H�N�U�'����/mZgv��gň_�4T���5���
����+ɰU��h��Qnsyk��nY�~��it��>r��=PQnsyk��n*w'_bN߈ݵYi�Qnsyk��n0���,0x�ݵYi�S��>�I2x�v�=�HC"zQ��� ԫ}/^�"�dI�?��ڸ�fb�%���mV��B�.�Xz$)�����>b�%���mVc�oK�SK��>������b�%���mVݾ!-��<7�;Fн�b�%���mV�N�Ƴ�tO�4b�%���mV`��(D�tO�4b�%���mVޞ����V�:_m=���p�"�2�SV��v������D�Oȝ����80D��6#�+k��	���r=�Y��r����&6ɽ�*<eɽ�*<eɽ�*<e!����M�h�L�E�6ω�*ܹg9�,�WM�4��BK_0Q����o=�����bC�x���b��6�-4�)�_π�e��A/�H87�]����H9������yõ�������x�r%=YF��)�xoĪ��㟰��TM�B"�O2�ia�s�a,4���?wƚ�����L��q���:v+5�S�����-���{Y\iqS��c�P/��+�ͼ�f���9TI��~-y7�����?�(<���Ef�]�k��-inh\�kܥ��q[��ղ�fǇz��X3������3e�X�Bh�W.����T�3@�ࣨSҝ[��R鯞�U�&4�h^�!������))�¼�H�4��l�ʶ���u�[��G1~l��҆2�1D���ɽ�*<eY[v�_�<��9��0#��J�= ȉ��f���9�)�]�찴�}0�@Z���ŗ AM��jt)�rj��+c�h
�K=4x�\�u+�n�/�G���q�����E�)��d��-QJ�ɏu��7)��S���+���M9�/"���S@�ࣨS,4���?wɽ�*<e�0�i�X�\$��I8�D��ݹ�V\_*X�#~v'�w�֬���AV�n��{M)����k����B ɽ�*<e�����d��1�d.�2���\&�k�I9^�ï�Lz�����K�P ��謋:���ڎX��S�2p[�������Ɯ�h�[�Z�~�qm�vo3�`ٮ��Z3{�~�g2H� �d�'x���S�+d��Ję���|��O��-���D���}�2���Y�����{������k��.���)Va&	3�W���%�THM�.���)Vw\��<���H��̞�.���)V$�os�7����-�B�j�^9}tq�",1�d��-QJB�j�^9Z�B[���Gk]91Ŗ��.���)Ve�V��u=oX�H�Nn?)���i�؁��ugň_����E������JZO<�
����+��
���WϓF���0�Y�~��it�û=55F���0�*w'_bN߈�
���WϓF���0�0���,0x��
���Wϓ��rP����x�v�=x�/φCi��۸Pp�%QB�2ƍ�zCr�6���	i�طt�"���l�w�a0�u,.姎��a���h
�K=4ɽ�*<eɽ�*<eɽ�*<e6��/�нf���10
����3,����;��	Զ����Qݓ˟s4�)�_π ����������'�e����ǄU���B(�{hԡj���	P�T����)���KS�$����sbRIꐦO�j$W.����|c� k�k��L�����`w�	�6�cx�\�uJ�fMw~�(�߷G�ey�q�ɚ G�Z[��� |2w�e�Q��kC����^��N2�{�&�����ڧ�ᦲc�����n��rɽ�*<e�m=����9қ�u;`J�d��-QJ��{Y\iq���Lt�c�/��+�ͼ�f���9TI���.�NH�����?�(<����t5��;��̲�E6�#
%��+��@�v;�z���v������D�Oȝ��QL�~Pw�	�6�cɽ�*<e'a���ˑ�#+�m�� �^[V�Cg�)�rj��+c�m<>�m�^�v2}&�PZ�n.{{�^��&��ᦲc�ɽ�*<eNM{9q���`���{�"M��
�/"���S�|����/�]�찴�}0�@Z���ŗ|ptjy��U��&�}�h
�K=4x�\�u+�n�/�G��`K�f���6��o��МB\'��ɏu��7)��S�Y�Y�����N�y��^C۪�Ml��,4���?wɽ�*<e&9��? ��9q:Xx3���^������eX�3%7|P���ޤ�]�찴�}0�@Z���ŗb��i���sX!�	�u>�o��P���� /"|�"�~���G>y�[]��ɺ��L]=�����6����_Ĳ�w�P � ��jY�q���36.^�d��%YC^2����ߐuX�q�0&�r�2����-���D�ߐuX�q�Dy秤_����RG�:O�ߐuX�q�$�s~e	Ӽ�j�<�U�q}���5�lv�G�0���j&��1��}���5�l��D�.��J ��u���ߐuX�q�RDk�,$�	��-���D�~�g2H� �c��Q�S������k�d��Ję��Jߌ���%�THM�%�G��ن������H��̞d��JęXq�!x�^����-��%�G���%`���yʏd��-QJ�%�G���\
|J:�Gk]91Ŗ��8����g�����6��o������@���쀏D�b+f���H�����+�J^�Q��	�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��,r�/�MeN�q�Xߣ�k �y����L�>��2��`χ�a$����^�M�"�ds��R��6G�2���-l	*v��I�,��؅��U>ɺ���V���/�#
%��+��Y��2�K+��+ v���Sd�~�fT�[V�`���S�)n%�\U�>:�NM{9q���\~C����jN�̓��)�rj��+cX��~?�W#��Jnj��?�{�/z�p�^(]e��#J�����`..
A���Y[v�_�W���P�#��6*+�'��^Ii6Q�v���%�;K�Raz�kC����^��N2�{�&�����ڧAv�'�B����n��rɽ�*<e���$�*�0.�#�d�!I�2dE�0(|�:B�2ƍ�zCCz���U%8�����}�\U�>:��VJUT���y�=R)��}�����\$��I8�����P�\_*X�#~v'�w�֬��������NJ��� ..
A���ɽ�*<e����옝�K��@��@��U��&�}�m<>�m�^�v2}&�PZ�n.{{3VUv�b�Av�'�Bɽ�*<eNM{9q��!�T9�k����S��N�y��^C���w�]�찴�}0�@Z���ŗ�mV�nzI�-�k�L�q�e���x�\�u+�n�/�G�YN�F�N�ꈍHg�8�3�F�K2f]}v���^B%aj�l�t�v2}&�@B1Y-�q f�&��������r=9xϞ�(��<�uO�%�t$�!P�N�Ě̆$�>qg�\XQH����c��~/^�"�dI��sZ��w4�v�Ѽ��B�.�Xz�ϥ�l<�S�v�Ѽc�oK�SK��4ȹ�5�v�Ѽݾ!-��<���K�v�Ѽ�N�Ƴ�+ �0���v�Ѽ`��(D�+ �0���v�Ѽޞ����VǛ
}���V����Jj�|Ĳ)�48lZ��_�E�+��43nb>�����Ϡ�����|;�NF��׈�`�%�����\#�@�]mp���V�B$g�Brh�!**��NF��׈�T٫��#�Z[��� ]mp���+ ���=��v���%�]mp����kB�]$l����A�%�jF���l�ʶ���u�[���F|����B
pfo����H�R�g��1-P��V]��%�ɽ�*<eɽ�*<eɽ�*<e,4���?w�+�ږ�F�X��X�+�)�ڙ�c �_`�ͨ�O��'��P�n�/ͻ�:||hy�6"pUw����^���F洰�-_ɪ�
a��1D��7�#J.�5�!I�2yh�S
cP�q>��Z�.����W�X��<R|=-}��&�rS�h
�K=4�&�;!��l�����k��-inh����P�[��ղ�f������������3e�X�Bh�Wd��ٰ#sf��Iă�Aҝ[��R�H�*��h�A�5B�	��U��&�}X��~?�W#|m9T�g�R?�{�/z�p�^(]e��C�]�Nf��h+�0�Y[v�_��H��g澁��Ş��i8�����}�"C�g�����6��o�����+~���0���))��h
�K=4����n��rj9PՂ�{�#f̨�~����������-��ɏu��7)��S��֧��`X��f�f��Iă�A,4���?wɽ�*<e��_NN��\$��I8�\�kܥ��q\_*X�#~v'�w�֬��-��?H!3<�䴗�.�h+�0�ɽ�*<e�������]/߷�W6�v����zI�-�k��m<>�m�^�v2}&�PZ�n.{{~25!��`���}*.�ɽ�*<eNM{9q���ܡ�,�'�%=��CTZ� g�+�����ʠ��6�L�d�[s�	�4�ڟ�}�}�(�L+'�w�֬��_�1��Ø��8B`}�FW,P��/b&�'�}�����֩�*��x`E%�N��|d$o���7�3]N|�F�j�!f��=oX�H�N�U�'����/mZgv��gň_�4T���5���
����+ɰU��h��Qnsyk��nY�~��it��>r��=PQnsyk��n*w'_bN߈ݵYi�Qnsyk��n0���,0x�ݵYi�S��>�I2x�v�=�HC"zQ��� ԫ}/^�"�dI�?��ڸ�fb�%���mV��B�.�Xz$)�����>b�%���mVc�oK�SK��>������b�%���mVݾ!-��<7�;Fн�b�%���mV�N�Ƴ�tO�4b�%���mV`��(D�tO�4b�%���mVޞ����V�:_m=���p�"�2�SV��v������D�Oȝ��C�����6#�+k��	���r=�Y��r����&6ɽ�*<eɽ�*<eɽ�*<e!����M�h�L�E�6ω�*ܹg9�,�WM�4��BK_0Q����o=�����bC�x���b��6�-4�)�_π�e��A/�H87�]����H9������yõ�������x�r%=YF����S,��m��㟰��TM�B"�O2�ia�s�a,4���?wƚ�����L��q���:v+5�S�����-���{Y\iqd������/��+�ͼ�f���9TI��~-y7�����?�(<���Ef�]�k��-inh\�kܥ��q[��ղ�fǕpᓖC������3e�X�Bh�W.����T�3@�ࣨSҝ[��R鯞�U�&4�h^�!������))�¼�H�4��l�ʶ���u�[������/2�1D���ɽ�*<eY[v�_�<��9��0#��J�= ȉ��f���9�)�]�찴�}0�@Z���ŗZ������)�rj��+c�h
�K=4x�\�u+�n�/�G���q�����E�)��d��-QJ�ɏu��7)��S���tB�jr@�/"���S@�ࣨS,4���?wɽ�*<e�0�i�X�\$��I8�D��ݹ�V\_*X�#~v'�w�֬��n�r#�O1{M)����k����B ɽ�*<e�����d��1�d.�2���\&�k�I9^�ï�Lz�����K�P ��謋:���ڎX��S�2p[�������Ɯ�h�[�Z�~�qm�vo3�`ٮ��Z3{�~�g2H� �d�'x���S�+d��Ję���|��O��-���D���}�2���Y�����{������k��.���)Va&	3�W���%�THM�.���)Vw\��<���H��̞�.���)V$�os�7����-�B�j�^9}tq�",1�d��-QJB�j�^9Z�B[���Gk]91Ŗ��.���)Ve�V��u=oX�H�Nn?)���i�؁��ugň_����E������JZO<�
����+��
���WϓF���0�Y�~��it�û=55F���0�*w'_bN߈�
���WϓF���0�0���,0x��
���Wϓ��rP����x�v�=x�/φCi��۸Pp�%QB�2ƍ�zC1�Y��N�?i�طt�"���l�w�a0�u,.姎��a���h
�K=4ɽ�*<eɽ�*<eɽ�*<e6��/�нf���10
����3,����;��	Զ����Qݓ˟s4�)�_π ����������'�e����ǄU���B(�{hԡj���	P�T����)���KS�$����sb�
T����$W.����|c� k�k��L�����`w�	�6�cx�\�uJ�fMw~�(�߷G�ey�q�ɚ G�Z[��� �/�ӄi�4�kC����^��N2�{�&�����ڧ�ᦲc�����n��rɽ�*<e�m=����9қ�u;`J�d��-QJ��{Y\iq�f��/��+�ͼ�f���9TI���.�NH�����?�(<����t5��;��̲�E6�#
%��+��@�v;�z���v������D�Oȝ2:(�@Հw�	�6�cɽ�*<e'a���ˑ�#+�m�� �^[V�Cg�)�rj��+c�m<>�m�^�v2}&�PZ�n.{{)���g~�ᦲc�ɽ�*<eNM{9q���`���{�"M��
�/"���S�|����/�]�찴�}0�@Z���ŗ��qy�6�U��&�}�h
�K=4x�\�u+�n�/�G��`K�f���6��o��МB\'��ɏu��7)��S���\`d����N�y��^C۪�Ml��,4���?wɽ�*<e&9��? ��9q:Xx3���^������eX�3%7|P���ޤ�]�찴�}0�@Z���ŗb��i���sX!�	�u>�o��P���� /"|�"�~���G>y�[]��ɺ��L]=�����6����_Ĳ�w�P � ��jY�q���36.^�d��%YC^2����ߐuX�q�0&�r�2����-���D�ߐuX�q�Dy秤_����RG�:O�ߐuX�q�$�s~e	Ӽ�j�<�U�q}���5�lv�G�0���j&��1��}���5�l��D�.��J ��u���ߐuX�q�RDk�,$�	��-���D�~�g2H� �c��Q�S������k�d��Ję��Jߌ���%�THM�%�G��ن������H��̞d��JęXq�!x�^����-��%�G���%`���yʏd��-QJ�%�G���\
|J:�Gk]91Ŗ��8����g�����6��o������%��:��쀏D�b+f���H�����+�J^�Q��	�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��,r�/�MeN�q�Xߣ�k �y����L�>��2��`χ�a$����^�M�"�ds��R��6G�2���-l	*v��I�,��؅��U>ɺ���V���/�#
%��+��Y��2�K+;	��7�8�Sd�~�fT�[V�`���S�)n%�\U�>:�NM{9q���\~C����jN�̓��)�rj��+cX��~?�W#�`���$��?�{�/z�p�^(]e��#J�����`..
A���Y[v�_�W���P�#��6*+�'��^Ii6Q�v���%���?��B��kC����^��N2�{�&�����ڧAv�'�B����n��rɽ�*<e���$�*�0.�#�d�!I�2dE�0(|�:B�2ƍ�zC�{l��E�_8�����}�\U�>:��VJUT���y�=R)��}�����\$��I8�����P�\_*X�#~v'�w�֬��+!�R��CYNJ��� ..
A���ɽ�*<e����옝�K��@��@��U��&�}�m<>�m�^�v2}&�PZ�n.{{��;���Av�'�Bɽ�*<eNM{9q��!�T9�k����S��N�y��^C���w�]�찴�}0�@Z���ŗ�)��.��zI�-�k�L�q�e���x�\�u+�n�/�G�YN�F�N�ꈍHg�8�3�F�K2f]}v���^B%aj�l�t�v2}&�@B1Y-�q f�&��������r=9xϞ�(��<�uO�%�t$�!P�N�Ě̆$�>qg�\XQH����c��~/^�"�dI��sZ��w4�v�Ѽ��B�.�Xz�ϥ�l<�S�v�Ѽc�oK�SK��4ȹ�5�v�Ѽݾ!-��<���K�v�Ѽ�N�Ƴ�+ �0���v�Ѽ`��(D�+ �0���v�Ѽޞ����VǛ
}���V����Jj�|Ĳ)�48lZ��_�E�+��43nb>�����Ϡ�����|;�NF��׈�`�%�����\#�@�]mp���V�B$g�Brh�!**��NF��׈�T٫��#�Z[��� ]mp���+ ���=��v���%�]mp����kB�]$l����A�%�jF���l�ʶ���u�[����C��A���B
pfo����H�R�g��1-P��V]��%�ɽ�*<eɽ�*<eɽ�*<e,4���?w�+�ږ�F�X��X�+�)�ڙ�c �_`�ͨ�O��'��P�n�/ͻ�:||hy�6"pUw����^���F洰�-_ɪ�
a��1D��7�#J.�5�!I�2yh�S
cP�C�6�vm����W�X��<R|=-}��&�rS�h
�K=4�&�;!��l�����k��-inh����P�[��ղ�f� �D�O�h>�����3e�X�Bh�Wd��ٰ#sf��Iă�Aҝ[��R�H�*��h�A�5B�	��U��&�}X��~?�W#m��3+� �?�{�/z�p�^(]e��C�]�Nf��h+�0�Y[v�_��H��g澁��Ş��i8�����}�"C�g�����6��o����~�#�y�Ip��))��h
�K=4����n��rj9PՂ�{�#f̨�~����������-��ɏu��7)��S����k3��f�f��Iă�A,4���?wɽ�*<e��_NN��\$��I8�\�kܥ��q\_*X�#~v'�w�֬���D;�k�<�䴗�.�h+�0�ɽ�*<e�������]/߷�W6�v����zI�-�k��m<>�m�^�v2}&�PZ�n.{{�t�3�2����}*.�ɽ�*<eNM{9q���ܡ�,�'�%=��CTZ� g�+�����ʠ��6�L�d�[s�	�4�ڟ�}�}�(�L+'�w�֬��_�1��Ø��8B`}�FW,P��/b&�'�}�����֩�*��x`E%�N��|d$o���7�3]N|�F�j�!f��=oX�H�N�U�'����/mZgv��gň_�4T���5���
����+ɰU��h��Qnsyk��nY�~��it��>r��=PQnsyk��n*w'_bN߈ݵYi�Qnsyk��n0���,0x�ݵYi�S��>�I2x�v�=�HC"zQ��� ԫ}/^�"�dI�?��ڸ�fb�%���mV��B�.�Xz$)�����>b�%���mVc�oK�SK��>������b�%���mVݾ!-��<7�;Fн�b�%���mV�N�Ƴ�tO�4b�%���mV`��(D�tO�4b�%���mVޞ����V�:_m=���p�"�2�SV��v���@�/�����R�)���6#�+k��	���r=�Y��r����&6ɽ�*<eɽ�*<eɽ�*<e!����M�h�L�E�6ω�*ܹg9�,�WM�4��BK_0Q����o=�����bC�x���b��6�-4�)�_π�e��A/�H87�]����H9������yõ�������v���y�1�$W.����|c� k�k��L�����`w�	�6�c,4���?wƚ�����L��q���:v+5�S�����-�1��zfA�kC����^��N2�{�&�����ڧ�ᦲc��VJUT���?�(<���Ef�]�k��-inh\�kܥ��q[��ղ�f���;��Y�/��+�ͼ�f���9TI���.�NH�h
�K=4ҝ[��R鯞�U�&4�h^�!������))�¼�H�4��l�ʶ���u�[����֙2Lx2�1D���ɽ�*<eY[v�_�<��9��0#��J�= ȉ��f���9�)�]�찴�}0�@Z���ŗ��ݐ�1)�rj��+c�h
�K=4x�\�u+�n�/�G���q�����E�)��d��-QJ�ɏu��7)��S��H!��/"���S@�ࣨS,4���?wɽ�*<e�0�i�X�\$��I8�D��ݹ�V\_*X�#~v'�w�֬�Ț�/�� ��{M)����k����B ɽ�*<e�����d��1�d.�bF�퉭�A��mt�[�t�r�'Q'9��O
W3���^������eX�3%7|P���ޤ�]�찴�}0�@Z���ŗb��iP�z,�JHy.��ׄ|�-�%�>����AKw�2�M�C���u���ДVkr����4\��]�찴�}0�@Z���ŗ�r��En�1�d�Ĉc�\��R*��\ؐ�V����d�ҹ[&���[��
����?�3�jb�&��B7YE}^�����D�h�|,G�N����FN菛�X��Q&fmt�*���	��Z��w�<Z���yt���#��W�}ѤD����8�3�F�K2f]}v���^B%aj�l�t�v2}&�@B1Y-�q f�&��������ᛵ���!z��/l�au��;����I����n�F�{FWS%�~�ǩ��[]��ɺ�lo�i�n@��vb!��wF�Q�k��/�v���������-[��,e/��S��R#l�{x����
j������k���gp��E�O�B�]t�$�m^�]|F	�N�"-w��-9c6p*���+�NG�Y�~��itQ��4'����ᛵ���K;.z���y{�ЯU�$Ņth���ĥ9���=lu��e�O+`��(Dr���4GH�]}i��%�~�ǩ���;7J���Xi!��߭vb!��wF�Q�k��/�RDk�,$�	��-���D�,e/��S��R#l�9`�G����^0�Phf��;ց����O�B�]tłr'����
����+ɩ��*[���9c6p*w�7TW��]���z�-$�������ᛵ����$����N�Ƴ̧th���ĥ9���=l�h�T<�&�������Ԑ�RBB���]}i��@�rj\�!.�kB�]$lX\AqQ����䢅L�����1VRKD�vQFƚ��������l�w���{A;�0
*�Ϝ&1�xAY{�#w�)3��Z������D���lkGpC��Y���U���B(�{hԡj���	[���F��sʶ��6L�h�UU��xr�^�i��zW-;�+j8ҝ[��R�?�mP_* >[����yB�VT�́����@��gpSPJeX.y$��#��?�(<���Ef�]��V�mB���x��{�&�|�D��U��&�}(B�W��ɽ�*<e�0�i�X�2���A`��Cr���]�BF'�̨�������n��rj9PՂ�{�#f̨�~���Җ LF�zN�����j9PՂ�{5���Y[v�_�W���P�ұ�Y:�f~w�)3��Z�������w�%s��l�0��NM{9q��!�T9���]'t�:.H.�4��(������S�,���МB\'�ҝ[��R�4r�k�\��4��{���
�S�E�y�݋�y�_(вy�B|�p�n����g��H8�������oCP�ٶ~xFB��;���K�Ѫ���HN�pu?�*i_�V/AY�X�@��Bi�Xƻ�2����"�+�I��A�x7����x�~��r G��ӌ�s���4�F4�t�eO��y� ��@�(|�˟QIB9/�I�\_tv�f&P�މl�p~rև]k<�E�I�.d����=(@���&?Vwn\�?�}ܴ�7'�PF(|ʮE��Ӯ�)��/�欿���<�N���4B���<�%�;['��ڀ�fh��n�4�ۉ�-.k���j�*Rq(/á���(��<��qy����~z``|YN�M��"%#k��-�[�6U]��$]���}~6�eW�^�Ԯ��%��o�a�U5)aF��WUw����x�Q�v{�-��N-�'��\c��Mݤ�Q�g�Ɋ2odq��3���
��?���� �A�����n uA�6[���n&?{<�0V+�+��~[�(��4Q�밈\f2lT�q�0N����<��N���h�-��MJє�Q�α,Ɯ�<�-	�30�5]ox��zs@]R/R�`�޷�'��4��^��M�)�qfy4_�I��u\״:�i\��DF jl�v���Weh�����O��L$���8����Q,d�P�Ӈ�>>���18��!�a��&�'1�C�eO��y� �
jR(�,s9�����4�R#l�X��2��s�bb�՞0WB|tn&K��!�
ځӏO�u�����K�~�6�ӑC#��6�\xO�հ���5�� �/j��_��2J���p��1�j>���p0�hi��j�h��4�ۋeN�b�v�w��b�	a��J�K� 6e�!/��bs� ��#&2Bna�&�Z��Ov� ���Ҡ�;��NE���w.�KL�k���IT��1�&����hx4�.�2w�C����p~rևb?@m̳�x�t�e-GT�)�q4X,�,�j48���ԙ���5�H�Q$�3��Xp���l��)c��&pW�,���A�����4��[C-�b2F����=_����������p0�hi��j�h��4�ۋeN�b�v�w��b�	a��J�K� 6e�!/��bs� ��#&2Bna�&�Z��Ov� ���Ҡ�;��NE���w.�KL�k���IT��1�&����hx4�.�2w�C����p~rևb?@m̳�x�t�e-GT�)�q4X,�,�j48��;�v����Q�����h�-��MJє�Q�α,Ɯ�<�-	�30�5M�
-JB�!�Ɯ<�O@�`�޷�'��4��^��M�)�qfy4_�I��u\״:�i\��DF jl�v���Weh�����O��L$���8����Q,d�P�Ӈ�>>���18��!�a��&�'1�C�eO��y� �
jR(�,s9�����4�R#l�X��2��s�bb�՞0WB|tn&K��!�
ځ��s^ 5$☼F&��U�~�6�ӑC#��6�\xO�հ���5�� �/F8���$���o Z\�9pKqfy4_�I9j�I)�N�~`�|�<�lz/�[t� H*�c�p��9�&�d³�Hެ�>����
��?���/i|�삫*��6��� uA�6[���� t�fXz Bۮ0� ���+�E������4��#�l*,���!�����p��M�HݹR'ť��l�W���_��ߧo�*�"���:���������l�z�=iv��&�Z �ʫ����Q#5 ���+Fo���	Ĝ�ա-<0;��~��I���4��^��M�)�qfy4_�I��u\״:�i\��DF jl�v���Weh�����O��L$���8����Q,d�P�Ӈ�>>���18��!�a��&�'1�C�eO��y� �
jR(�,s9�����4�R#l�X��2��s�bb�՞0WB|tn&K��!�
ځF}7��h���RV@7���Xp���l��)c��&pW�,���A�����4��}�
��9"w̭��#/D^PtH)�|/L�$ɠ_M�x�蹹�Hl#[ė���D�h���\�����eO��y� ��W-sD'�4tꦘ���R#l���w�%�<&qj�Iؾ��$s:������8��^R�������߳�_ەU�6����7
�E�Yؽ�&�b!B����Ż�5"rb�=�[Z��� �1��:��h�-��MJє�Q�α,Ɯ�<�-	�30�5����-�NCGk]91Ŗ��ad�֙��;V�l�Un�f�i��OIu9؎w_eC������4x{�B<+-T2N_PzB �k�3W��1�&���N�9����?��1t�p~rև-��䇧wbZ�vH�fs{�̦I�_���
�C���K��X�qǑ5�X�Yg�W���NN3V,q�̡h��q5��x�٩Q�6��r$LZ{�m0�m�����j�C�
]�� �!k��B�,����
�D�:&#��51u�څ��L�I6�ތ`����)F���ƋY-(1��
17IEV�]�ҍ��r�M����chaW�T%�)��O?�Y+�IS�a�?S�]������ˢ�J�� ��@�)�_tR��Xw	r�j�5��B���bs� ��#gc���_v!��N>l��a{�0�^'�S�V��|�?�>�P�S����0_����j�$�7�����j�C�
]�� �!k��B�,����
�D�:&#��B�.�Xz2J���p�'��b��M��"%#k��-�[�6U]��$]���}~6�eW�^�Ԯ��%��o�a�U5)aF��WUw����x�Q�v{�-��N-�'��\c��Mݤ�Q�g�Ɋ2odq��3���
��?���� �A�����n uA�6[���n&?{<�0V+�+��~[�(��4Q��ݪ6�E�=`!m����Q�����h�-��MJє�Q�α,Ɯ�<�-	�30�52�r�nPq|F	�N�����!�cqfy4_�I9j�I)�N�~`�|�<�lz/�[t� H*�c�p��9�&�d³�Hެ�>����
��?���/i|�삫*��6��� uA�6[���� t�fXz Bۮ0� ���+�E������4��#�l*,���!�����p��M�HݹR'ť��l�W���_��ߧo�*�"��2���������7PƏRP��Fǫ�%�t^n��y~��	s��cU�K����@��Y�~��it��e�J,�Iތ`����)F���ƋY-(1��
17IEV�]�ҍ��r�M����chaW�T%�)��O?�Y+�IS�a�?S�]������ˢ�J�� ��@�)�_tR��Xw	r�j�5��B���bs� ��#gc���_v!��N>l��a{�0�^'�S�V��|�?�>�P�S����^2��$q�\6q3�]���v���!���dC���e��آ�e�M!N���f��mga��q���� T�M�|��<l-�+͘3+1/�s�<���U�P�o�P�[�omK@�Y���V$���`i���8V�����6~8� VQT�!��t̞�����a�}[�t9ƙ�]�?M=�R�i%���XǮ�O��L$��F*�T��'�]J0:���Z��C����?���k&X�L��iԴ�#��Pg�[�}BJg^���j�C�
]�� �!k��B�,����
�D�:&#`��(DG�BT6�̢;V�l�Un�f�i��OIu9؎w_eC������4x{�B<+-T2N_PzB �k�3W��1�&���N�9����?��1t�p~rև-��䇧wbZ�vH�fs{�̦I�_���
�C���K��X�qǑ5�X�Yg�W���NN3V,q�̡h��q5��x�٩Q�6�P(4 U����� �1��:��h�-��MJє�Q�α,Ɯ�<�-	�30�5+�&��aC��ۅ�{<d�Ly��.�#/D^PtH)�|/L�$ɠ_M�x�蹹�Hl#[ė���D�h���\�����eO��y� ��W-sD'�4tꦘ���R#l���w�%�<&qj�Iؾ��$s:������8��^R�������߳�_ەU�6����7
�E�Yؽ�&�b!B����Ż�5"rb���$F�nX�#��=G�[��#U)���Xp���l��)c��&pW�,��{i�������K�����k�I9^�ï�Lz�����K�P ��謋:���ڎX��S�wY���=�@Z���ŗG.|�w@����Ɯ�hZ҂=����u�[���z&Ƙ�����#ڄ�֐ s:_�OP��0��x�\�u^��
:�*�~�sh-���b}�����Q^�|�,Ksk���Z���-\dE,>������D\ȯ�?��N.̹��_<��D���&ZReX�NM{9q���w��ѹ����)��Yj�ԢqL�A)�rj��+c�h
�K=4����였m=����9�n��4�}��;#�l<�%K\�dջ�ZXd�"uUI�,-Я��`K�f�<������;q���aj2�1D���,4���?w9�C�)���J�= ȉ>|
ϒ���sm���	�AE
!�x�\�uH�*��h�Aa���d1�W�D6�fD�$�qh+�0�Y[v�_���]/߷�W6�v���������s$)�	�)��NM{9q�������i�����1�����S"�E�����yO]�&��I���R��A|`�$������kȡ�B,ŭ_
j�����ͬT$OeMS���s�C�罤�9.�f�i����
D��H7����{�ƥUuh��V�g5D�l��9q�X�:׮�5:��KL����z�>�4[���{u�^ק��}�{�ʘ��SD!��Ю���0�V�٦�����2���X�����wD`֡��y����"�m���F^��`���#H����^'�2����:W�0s�����S�_>gN�-�:'��$+���G(����^Le�0�[��z����jcbb_�B�,��y8f���B6Km���'�5uEq_�<|7.���|N;X�^�I�[\o|�o�����|"ÝW}�utiO����+�%�Q)=d���E,��h��DZ�x���F\��w�0��8w���c�Y�l�%�tB�*��� �&&s�:v3�9?k����Q������L�����p�N_�qe�
��>̊��%�
�T���k���g���*�F/��q+�\��$|?G��a�G�x�D�9ϑm�eQ���9*Q����� P�7+��$-���G[�z�A��ie�\#�_Hc����'d����uC)�E���Q�0)Dm*
kma��ݑ�`��N��X5/�)I�|��o9�H[��UF�n]h�^�o��p����=����+P
���(�5;B�W��M��v��E�`�w$�P��j�:�mheˣ��:��?Dg,2ms����{Ue#T&�ީ�q�� B����ĸ��Y������kȡ�B,ŭ_
j�����ͬT$OeMS���s�C�罤�9聯�v!�������k{��Ty}�zj�"��0��U��j )���.s���2D��%_�y��N�[\��NT��>n.r�P�S��И]h����,��D�se��L���Ӡ��B:l��9q؟��?��6\F�߉�}3z�s"�!6���f����!Lؒ&�bL�.��. ����lB��,zyj���0_��A�\��B�N��%졖*��j)?��(a�����@��$�G#�ӵI�0��#Ҟ�s�-I@>������BP�\_�0'���I"ʈ�W�rB�������i0aXK��2��H����D���i�6 ��Z�)a��\ `L����B)JǴ��	ĭ��n�W���\?�R�?3�h0)�E�Z��(w
�7`�	�6�����C��F���Y��U��>��M���2�أ���Q������L�����p�N_�qe�
��>̊��%�
�T���k���g���*�F/��q+�\��$|?G��a�G�x�D�9ϑm�eQ���9*Q����� P�7+��$-���G[�z�A��ie�\#�_Hc����'d����uC)�E���Q�0)Dm*
kma���t�jp�]$u�	8'��v�eMV�z�U܉����4�=z��F		DAu��6YhzoC-x�i���
V�r&A�V�6�.j���|R��Ǥ_�|�P��L���Xj��)�*��e/6�5��0�Lu.���v�� �H��{2��ħ$(�MZ��Qa-u��B���0���-��nQf�z]�R鮎����|�Z����z%u=���a�ҡ����U�포�	W����~�	��>�d����_�|�a�*��J=�u�Jm�X���F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8� |ݰ&���_>וL�>w�@g��:dU��9���o]�5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�/I�T���cψ5���4ݾ��䐐��F���VF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�LB�X���`,ȩq/]������˫'mdO0?Y���W<:K+>[����/�p+�3���^������eX�3%7|P���ޤ�]�찴�}0�@Z���ŗc,�*
:�PZ�n.{{b��i��<�a�]�;���	���V=�"�ɽ�*<e���=s� HK����6�͟^O@����c���&��@��Z�ݐ;��?t����/s!_ǁ�3�A;Q&{���s�-<�������8�Cl#�8H�rpl��g��#��b��s��Α9��������[Tװ����yK80�L^ʔ��.�"3$��>����Y7�:f��$E�Ylka/ځdm�İ����O�Rgo4G+jvϥ\�k$b ��K�Z9"^�iW?54�wi'��/�Ns�48&����E�Ylka/ځdm�İ����hR���8��S"y�B�L,��y�C3-j4�	y�G�Vgl�%��q����
>zby"�aJ��D����޼�\?�>�.��5������x�! f�SL��(�|�;�S/܀J���[���ު3�*�q�3m��x��\4��V�ɽ�*<e�wi'��5"�_ Nɽ�*<ed*�cHа^A7FO�JNY��s����p���+�	����Yo�P������F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8����DW�S�ph9!�4�hԚԾ3��Q���d�O��]��Ɩ<���l�ʶ���u�[���~{]�*��s76?b=��K�XLT>��:��B;ߐ��yם�A�<�Ʃ6��/W�����a3m����@����xw��E.8Ԙy�9ɽ�*<eƚ������=��c��v���K-�c�G+*�ü�L���1D����:ʉ$�Hl�&^D~����� ��#*ɽ�*<e]�P�.�Fx����Q������N���6����=�]�P�.�F� ���	/����N���r� ��v���ѫeFaȫһAm����N���Jvk�h\�S�Ƃ���dm�İ����:-j���Uj+����1�2P'L�E.8Ԙy�9ɽ�*<e���r�< ��ϫ)��;��t�^	�#�x0U�o\�I;���ɽ�*<e`ύ���#��̿u���E"��R:�����V�[�?tR7��&e���Fa<a��I�IT���/�_��I���� �8+׊����F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�ol&���rl��+����-_�5a���`�
�������F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8���n�.:�	~���`V�f�Bƚ������5���Awo��o�x����&���#����DH77j4�+�(�T	�]�P�.�F�sE��@���a�Iw��SCR'3C}�/��cF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^��J��m ����V�O	�k��i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S�j`▘9�E����_H2x���]L�E��2� �p?�G�^��A�Y��g���{
>zby"E^Ip������).��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e-� �FȤ��'�9�3���Ъ���=E��Rx����琘���yO]�&��I���R��A|`�$������kȡ�B,ŭ_
j�����ͬT$OeMS���s�C�罤�9.�f�i����
D��H7����{�ƥUuh��V�g5D�l��9q�X�:׮�5:��KL����z�>�4[���{u�^ק��}�{�ʘ��SD!��Ю���0�V�٦�����2���X�����wD`֡��y����"�m���F^��`���#H����^'�2����:W�0s�����S�_>gN�-�:'��$+���G(����^Le�0�[��z����jcbb_�B�,��y8f���B6Km���'�5uEq_�<|7.���|N;X�^�I�[\o|�o�����|"ÝW}�utiO����+�%�Q)=d���E,��h��DZ�x���F\��w�0��8w���c�Y�l�%�tB�*��� �&&s�:v3�9?k����Q������L�����p�N_�qe�
��>̊��%�
�T���k���g���*�F/��q+�\��$|?G��a�G�x�D�9ϑm�eQ���9*Q����� P�7+��$-���G[�z�A��ie�\#�_Hc����'d����uC)�E���Q�0)Dm*
kma��ݑ�`��N��X5/�)I�|��o9�H[��UF�n]h�^�o��p����=����+P
���(�5;B�W��M��v��E�`�w$�P��j�:�mheˣ��:��?Dg,2ms����{Ue#Ty� �I�quȯ����2���Ե+�ynB�;{�7�$$x<n���.�?g`k��fL7�x���{��I7�������j){Db�Ԫ�N�l$ku�,V z�C�_CeL�f�ZSl�Ȅ�{ڪ0��!�41ҕ�G�9����DC�#�/e�x�P�f��H�H�i�YEK�x7^LX�1�{��F2]�J8�F2]�J8�F2]�J8��<�2��M!�Q{L�������R�F�dH��su�~t�F��� T���ڭ�ݱ��֜,dY�,����սX/N�D���'�=�Uq+,�o��v��r��ԋ5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8��"�iS{/E�́7�׈�|�.��b=�D2�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S�X<��a5���I uA�6[����S�2͙gG�7W��d(�e��'_>g�Q]e8�3�F�K2f]}v���^B%,˛e1?�2g\ɳ���q f�&�,/�z/�X� %��N)O�yf�!ɽ�*<e~��\�/����S����t^����?�����t��&3h�t�U��"�W̌a�����Kx����(���ؙQɽ�*<eܞ��G��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�S<��1���F2]�J8�F2]�J8�F2]�J8�F2]�J8��<�2��M%mD*��+�G�O��d��[�u�aH��[�ї'�h02%Qk!F5ğ��ه�rݶU���e�y0ѷ��h���9kZ���v�t!cJ(�Z�0�W4iE�a�Q�e:���,�	z��$�P~F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8����Ѹ��:����oz)���ʠ��6�L�d�[s�	�4�ڟ��s���T� J�F�{��8B`}���^b�AaKC��ଡ଼�F2]�J8�F2]�J8�YZ͆ˎ�0�`��D�����F2]�J8�~�&T�S�5��Oh`M�p�+0�{	i+����w�~x'J�9��E�]�Ҽ�w	^�R�u���T+���-w�~x'D{�1��K��~��.�hjᔇZq�c]�Ҽ�w	��؋x�Hg��*KvcJ��KE��۳���F��a�sT7u��QӛE,�����@O�.�^<�
:�ɽ�*<eɽ�*<epH[��V�"�#F��87U*���g5��Oh`�wo�	h�[ɽ�*<eɽ�*<eh���|s�b���<���^�NI|	*�eF9YH,ɽ�*<eɽ�*<e!ՠ��s������V<�κ��_i�ܛ�|�F2]�J8�	C7��3�^�˽�c����vZ�R�C��ଡ଼�F2]�J8�F2]�J8�M��1�����f�[>���ɽ�*<eɽ�*<e�����`�v�<����M��1�����f�[>���	<�9��i��<f֩����Bo�� KЋ��7DG��n�jF��72L%hQQ����5���VL��8����c����������)D���u8��I�J���W<:K��{v���ɽ�*<eɽ�*<e�[7%�`G5�td'P�TT�I���W<:K��{v���ɽ�*<eɽ�*<ek�e�=M�����<���^�NI|	*\�I;���ɽ�*<eɽ�*<eɽ�*<e����t�dHL�`I\����N���6����=�ɽ�*<eɽ�*<ey��ٕf�#���k�L�����N����/Xb,k��T+���-��{�q�kI+�<r���H��8xyb3���D�u�w��5��M����Հ��-Ncź9�/�闺IOz��0�۳���F��a�sT7u��QӛE,��=̦`o����9��ɽ�*<eɽ�*<e�K,V[d}�g9�bV8��+ Z؋$��,!����9��ɽ�*<eɽ�*<e�K,V[d@h[�T��7U*���g5��Oh`�wo�	h�[ɽ�*<eɽ�*<e��S�c���x����Q��M��1�����f�[>���ɽ�*<eɽ�*<e�����`���x�Z��)M��1�����f�[>���	<�9��i��<f֩�}'{�P"E�� KЋ��7DG��n�jF��72L%hQQ����5���VL�o9�$�pD���������)D���u8��I�J���W<:K��{v���ɽ�*<eɽ�*<e�]�����MG5�td'P�TT�I���W<:K��{v���ɽ�*<eɽ�*<e�;<�]iT���<���^�NI|	*\�I;���ɽ�*<eɽ�*<eɽ�*<eQ?%�yIdHL�`I\����N���6����=�ɽ�*<eɽ�*<e�*B<W����k�L�����N����/Xb,k��T+���-B��aq��+�<r���H��8xyb3���D�u�w��5��M����Հ��-Ncź9�/���i���۳���F��a�sT7u��QӛE,��=̦`o����9��ɽ�*<eɽ�*<e�K,V[d�0*����V8��+ Z؋$��,!����9��ɽ�*<eɽ�*<e�K,V[d&Py�eH�7U*���g5��Oh`�wo�	h�[ɽ�*<eɽ�*<e�~��xӴ�x����Q��M��1�����f�[>���ɽ�*<eɽ�*<e�����`�a���~��M��1�����f�[>���	<�9��i��<f֩��	x-�� KЋ��7DG��n�jF��72L%hQQ����5���VL��{/U Qz����������)D���u8��I�J���W<:K��{v���ɽ�*<eɽ�*<e�BI�"�NG5�td'P�TT�I���W<:K��{v���ɽ�*<eɽ�*<eC�1B��m3���<���^�NI|	*\�I;���ɽ�*<eɽ�*<eɽ�*<em�%���dHL�`I\����N���6����=�ɽ�*<eɽ�*<e,ѥ+�����k�L�����N����/Xb,k��T+���-��d��F��+�<r���H��8xyb3���D�u�w��5��M����Հ��-Ncź9�/��Ԉƹ���۳���F��a�sT7u��QӛE,��=̦`o����9��ɽ�*<eɽ�*<e�K,V[d���!@%XrV8��+ Z؋$��,!����9��ɽ�*<eɽ�*<e�K,V[d2Ϭ%���7U*���g5��Oh`�wo�	h�[ɽ�*<eɽ�*<eS�?w5�$Xx����Q��M��1�����f�[>���ɽ�*<eɽ�*<e�����`�  H�L��M��1�����f�[>���	<�9��i��<f֩�� @��;��� KЋ��7DG��n�jF��72L%hQQ����5���VL�Kb�������������)D���u8��I�J���W<:K��{v���ɽ�*<eɽ�*<e�r�1�CZ�G5�td'P�TT�I���W<:K��{v���ɽ�*<eɽ�*<e���]��Wp���<���^�NI|	*\�I;���ɽ�*<eɽ�*<eɽ�*<e��� N�9dHL�`I\����N���6����=�ɽ�*<eɽ�*<e=��sL���k�L�����N����/Xb,k��T+���-�%�z�?+�<r���H��8xyb3���D�u�w��5��M����Հ��-Ncź9�/���De�Fi�۳���F��a�sT7u��QӛE,��=̦`o����9��ɽ�*<eɽ�*<e�K,V[d�jz��kWV8��+ Z؋$��,!����9��ɽ�*<eɽ�*<e�K,V[d�x`�Y7U*���g5��Oh`�wo�	h�[ɽ�*<eɽ�*<e�J�?Q�]x����Q��M��1�����f�[>���ɽ�*<eɽ�*<e�����`��l�����M��1�����f�[>���	<�9��i��<f֩�'m8���� KЋ��7DG��n�jF��72L%hQQ����5���VL���������������)D���u8��I�J���W<:K��{v���ɽ�*<eɽ�*<e�7��7G5�td'P�TT�I���W<:K��{v���ɽ�*<eɽ�*<e1�矉ʠ���<���^�NI|	*\�I;���ɽ�*<eɽ�*<eɽ�*<e������dHL�`I\����N���6����=�ɽ�*<eɽ�*<e��.;�7����k�L�����N����/Xb,k��T+���-�F��vr+�<r���H��8xyb3���D�u�w��5��M����Հ��-Ncź9�/��T�,�֗l�۳���F��a�sT7u��QӛE,��=̦`o����9��ɽ�*<eɽ�*<e�K,V[d�]T�� [V8��+ Z؋$��,!����9��ɽ�*<eɽ�*<e�K,V[d�Y�=`,	7U*���g5��Oh`�wo�	h�[ɽ�*<eɽ�*<e�����P"x����Q��M��1�����f�[>���ɽ�*<eɽ�*<e�����`�]R�z�.k؋$��,!����9��CCgm�0�v��x�\�  i�ĕe��J�)��KBaiUj)��}	�c�hk�����N���g��� ��}@'��ono��b���z�g�-L�����S�4(8��pMM��1�����f�[>���ɽ�*<eɽ�*<e�����`�U�V�]�$V8��+ Z؋$��,!����9��ɽ�*<eɽ�*<e�K,V[du��/�\�_��F���]�Ҽ�w	�B�a�h�ɽ�*<eɽ�*<e�����`��앫�;`pٞ8���72L%hQQ��p��u��dɽ�*<e�p\�Ì�~rW蜠�kG���R���Kn�:O`��y%m��^7������(
�C+�<r���H��8xyb3���D�u�w��5��M����Հ��-Ncź9�/���dkX�����u��ּ�>Gc���l����-$*�5����x72L%hQQ��p��u��dɽ�*<e�p\�Ì��(N�Ȟ��̸B����NI|	*�Kn�:Ou
����.ɽ�*<eɽ�*<e]��ޥ�K�am@�nh��@�;�5����_k`ɽ�*<eɽ�*<e�p\�Ì���s��q����!\�C��ଡ଼�F2]�J8�F2]�J8�YZ͆ˎ�C����ß)��t#s!��C��ଡ଼�F2]�J8�F2]�J8�z�����& �ێr-k!�ex��>h��:�R��@�ԧQ����3��y�<{��o?�N|B��`�y��ܳ���8�v`wQ�s2l�f��K9!0ޱ+]�Ҽ�w	��f�jd�p�x���z�k<'����	�����?r
�x�1;����yf4�H�+_8�,���3�d=�� �;�"�<�*ʣ�Pwf����XS���5��+@G��p��E�Ͳ�������B�s=c@�LT2-T��#b�t�U�bH��*�?�Vl��n3�@P��7.*��'�|m����/��A+L*i��<!����w�C��ଡ଼�F2]�J8�F2]�J8�YZ͆ˎ��<i$ ?C��ଡ଼�F2]�J8�F2]�J8����d��X��[��Ƹx���]L�E�����`�#
%��+�ɽ�*<e��v~���ö�#5�����`�8�� �a�ٰ���˫�
�;>��G5�td'-�f��ݬ�K,V[d"V��A|m#��U��Z����˃�6��Rb����������`��8����c�[��%�w/_���y��l�tt��h��xp-n��o8^N�DXɽ�*<e$�EC���j�<�U�q;��N+ށ��BSҧ��{� ��Q}!�Lڜ�e3q��Oɽ�*<eg��E{j��49�iv (;��N+ށO ��sye�ɽ�*<e5�ε�����̸B���#�3�$� N�s��<��G���"������p���P[�q�I��K�am@��I�)X6vZ�%�MO�^p=�ɽ�*<e��b]�����B�"���;��N+ށ��BSҧ��&p+��Q����[1�W�4�b�z�a�h�H?�..+`��r���4GHB9Hl�+s���=�k��x��KC�f�.:!��ʞ�4�b�z�a�{g!��{��!I�2r���4GH�n �u�HY͌r�����{g!��{������d<�2�>��1c�XO�_ag�̸B���ثK*3�ҒHw$�����"vЅ\��Y�5�8��,#D7��K�am@�p���b�!��{g!��{�,�o��vr���4GHB9Hl�+s��s�Gv�<���?���3�����t7��K,V[d�{�v�%tɽ�*<e�����g#!x%q�&N�f�r4� b���ʀ�c�\��K,V[di�{�r�Oɽ�*<e����O�. ����K,V[d�0*����V8��+ Z���������d<���J�ܰ�r�p\�Ì����(��mٰ���˫��bvz�*�"vЅ\�-�f��ݬ�K,V[de����G�c�т����,�o��v��D5��L����(*����p���*B<W��q]�iʳ1Q��K��T3�_��G�(�ݣ�L�C�NX�Jj�*��Iv3C<����p��!m`h�`���������Q��K���s~;fT����p���ǃ'v#h[�!�(I�{�0�p ���؊��SV8��+ ZA�Y��gC�1B��m3���<���^Ƽ�A \�������^���"������p��%���ZdJ�J=���Q��K��T3�_��G��zwle7j��t�U�l�I�J����֗� q����P���*��cJ��KE��d	@���n3[����8(^:��>�PRL㥡�S�?w5�$XY��# N����*�����KT���V�)iS�?w5�$X"�#F��8�⠡��RJ��c��!�(I켗���������`��<sEvT�����of��Z�91�����<���^ثK*3�ҒS�?w5�$X��K�`��*��cJ��KE��*�Wji��������q��k�K�p\�Ì��'��pD	�Nd"�O���bvz�*��K�` M_�-p:'�09k� �`����?Ԥp\�Ì�� @��;��ɽ�*<e�bvz�*8�d�	���p\�Ì��zH�8��m�B���?����V"�#F��8O�^p=�ɽ�*<e���7��w�V8��+ Z;��N+ށ|M��t+c��J�ܰ�r�p\�Ì�������;��X����bvz�*��K�`�d�����A����^�ߔG�=�� 6vt�uצ���-����ؖ��u F�yz�G��EF��k$J�]���:�ߔG�=��xw=�+B��b��M&���ؖ��;�Y��##A�Y��g�C-w:��G5�td'QZv�i��`MlZp
T�m�B���p���b�!�X/���gD˃�6��Rb�SFt�a�r�=_V8��+ ZA�Y��g���9_V��Jd�q/ݼ��ؖ��u F�y�>�׭���ϒ0�-�m

c ������`��9��{�} ɽ�*<e_���y��l:E�D��zi���C?+�.\2���0��k������`���:���ɽ�*<e��v~���ö�#5�����`���pC��v_ٰ���˫�
�;>��G5�td'-�f��ݬ�K,V[d�-4���z�#��U��Z����˃�6��Rb����������`������[��%�w/_���y��l�tt��h��xp-n��o8^N�DXɽ�*<e�e�l�0���j�<�U�q;��N+ށ��BSҧ�6ͼޑ|��}!�LڜIX��\@ɽ�*<e�����mà49�iv (;��N+ށO ��sye�ɽ�*<e[,]!u�K;�̸B���#�3�$� N�s��<��G���"������p��P�4fR��K�am@��I�)X6vZ�%�MO�^p=�ɽ�*<eT`�*!�z�B�"���;��N+ށ��BSҧ��&p+��Q����[1�W�4�b�z�air{�:d�..+`��r���4GHB9Hl�+s��ޜ�w��8�x��KC�fK�ʤ���p�4�b�z�a����FXY��# N����*�����KT���V�)i��S�c���8�� �a�ٰ���˫�
�;>��G5�td'-�f��ݬ�K,V[du��/�\�_ٰ���˫��bvz�*�"vЅ\�-�f��ݬ�K,V[dR��{�F����X����bvz�*��K�`�d�����A����^�ߔG�=��,�k0=/..+`��r���4GHB9Hl�+s�1Lk�n�7�n3[����8}C�q(�1H ܷD�҄�����`��g�I��ɽ�*<e����O�. ����K,V[dO�3��qwm�B���?����V"�#F��8O�^p=�ɽ�*<e]��ޥ�K�am@��I�)X6vZ�%�MO�^p=�ɽ�*<eEgV����J�J=���Q��K��T3�_��G��zwle7j��t�U�l�I�J���S�c���!!,b� 2ɽ�*<e_���y��l���2[��i��iX� b���m�ǐc8�v��,��-��KC�F2]�J8�F2]�J8��� �z F7W�[j?��&�n!��*�D��|F2]�J8�F2]�J8��a��T�лV�|�®��o\ע�Q�嘄�^旿�]���L �ց�5��X���S~Ti�i��/�e/W�y�\���'{�5r{�
���ji�+L*i��<�<�C�X���+g�6��Wm*�����Q� �p��#@\0HM�(���퉢\DԷ��J}��Pj]��w��\�Y��߼8��2�% K�>Ѻ٤tF�(�[�v��6��D�SG1�KW�%b�MW�樳T�2+��@��^/aÊ,���kޝ�n?�����2����¡����V�}����u�9ݓN�O���-^T��.Z���Z��Fs�5t����?5лV�|�®��o\ע���ާx�t|z#�*C�M1�L �ց�5��X���S~Ti�i[/�uF_��F��,����'{�5r{�
���ji�+L*i��<q��4!��_Yw��uZ_>Ѻ٤tF�(�[�v��6��D�SGYi����=P�t�)Z��vt8�@�Jk�N*�%����u��_a������(yN�!���BSҧ�{j�З\�O���-^T���z(k�En������Uj�5�h���spoz�X�}��R��Z�J���F�c�q9r�T�?:�;���A��#�P:\����u)�QX^�2���@i"M6f��������5��	"	���?��o��N�1�a�g��ۓyP������1��
O?�p٫j��"�yL�x���Ys�}�q��?Xٵ��5�,����F]�J�������	UQQ*rb�5��6��uF�p�	_�P塙@:/!M_[V�I'�
n� 70^�d�e»�-0^��,�:�	S�uP�M�zK!�g٪�'�)��F�p�	_ى�#�9�$�oWU� ����L�m�C��#��;����B�	?�gwC�N�O�lK���K)��F��P������_#Ǚ��R�����'c.�	?0-� ����Jv���,����@p~�@oH��{T��qɮ����D���,%GJ�=�rW�K�v��|�5������zWG����ʙD�0@]�����>'�6�*�q�t������ϩU�R�4�t������:Wp<!���I��d�>�r=D�9�)�Ί#|�Ӏm��!Q	s>R=��@�wG�ɽ�&���[�O�VG/"���@V��"W���à\j����f���ԝh<K��}|�?�M��\%i�������E�!��o�8���RX<���O��"P)�6�m�`�� P����Y6Z����*y����,��/�&�5K}�*���ՙ��e'�������s�SŠ��z��Qd_No���?�%6=����e���w���t� �l�I/Ό%��c�q9r�T�?:�;���A��#�P:\����u)�QX^�2���@i�I/Ό%��c�q9���I|�� �V� �s�'�4s�����2s����	k��;l��O����S��mCSfe�%T00�ѐ�ͤ���]����%ޮ+x�(+M%Y�f"h�ۓyP�� m���� Դ��[��Os�w�F��֕pR�Lʉ/[¶���`���c��� �	[�w:���ע��������t��E�̎����D�<L}ڈ�����dn'y&���3��ͨL���K��a9q;���]��e�G<���ߤ#����ө�((|�w��M{� C<�ls���|����䋇�æ��tg������a��4W%��g���$�-�����Mv�'��X�)����qӬ�\ԗ������nx�I��	n�=��ϝ�p:�ɻtpe��IO҅�QҔ�n�zWG����ʙD�0@]�����>'�6�*�q�t������ϩU�R�4�t������:Wp<!���I��d�>�r=D�9�)�Ί#|�Ӏm��!Q	s>R=��@�wG�ɽ�&���[�O�VG/"���@V��"W���à\j����f���ԝh<Kaչ�z�Mf%�l�J�����7N?aJC��B���ڡ��n]h�^�o��p����=����+P
���(�5;B�W��M��v��E�`�w$�P��j�:�mheˣ��:��?Dg,2ms����{Ue#Ty� �I�quȯ����2���Ե+�ynB�;{�7�$$x<n���.�?g�} <Pr=~��>ҀVh�.v�#?kS�x���{�1�	"�Xߊ��l.m\5 �Β����ܔ������^u�{�=.��x�bW� ��:���ƺ#�FE��7�R�b=�D2�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S�?%6g?��ӣǠ>�Q�7�K��7X�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�/I�T���cψ5����4���m.o}��y��X�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�S(W�!������R����V��j	>Yn|��o6�5��M���� ��Ftɽ�*<ek�I9^�ï�Lz�����K�P ��謋:؆(�Y��b��i��<�a�]����\�p�i[�Eg�+,ɽ�*<eM��h'��˥�(��ZW�wucV�8ł�� �/_d"['�M��UEN,�~�v��� l/�M��HH���!��1vHt�!9@�73qF�[��0�ZM��h'T6����1�'�4�&�j�+�.S�℧��(��*�D8����,���3�K�ٷz_����Z���`?�8+.
�@�ɽ�*<e�Go�ҁ�h� K��3������8a�-_��f�xr>����C�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S��8�:o��k�I9^�ï�Lz�����K�P ��謋:؆(�Y��b��i��<�a�]����.�g{kX�1�{��F2]�J8�~�&T�S��!��(�V���6-������F2]�J8�F2]�J8��o���ٽ�5����_k`ɽ�*<eɽ�*<eX�����M � ���	/5��Oh`)���Q����v��x�\����.�ȅ�J�_���G�P�!R����R�7uh��F3'���]�Ҽ�w	�B�a�h�ɽ�*<eɽ�*<e�/(���iG5�td'P�TT�I��~��Wɽ�*<eɽ�*<e!ՠ��s|Gb��f	>��F���M��1����.�^<�
:�ɽ�*<eɽ�*<e7�'#GۭZ�׈y�WP-��KC�F2]�J8�F2]�J8�	C7��3�^�˽�c�Zء�خ'�5����fF2]�J8�F2]�J8�;Pj]p`ޫi�q�k�אɽ�*<eɽ�*<e>�t<sa�'���k�L�����N���	<�9��i��<f֩����K�=M��1����a�a�_��}@'��on���g�@PdheX��T��eF9YH,ɽ�*<eɽ�*<e[�Q�����d<�s��7Z�5��M��̠wo�	h�[ɽ�*<e�p\�Ì���W���7U*���g5��Oh`�wo�	h�[ɽ�*<eɽ�*<e4Wj̼�Шc�e[�J�5����fF2]�J8�F2]�J8�)V ٥�DkF�iZ���CA�0>��2*�D��|F2]�J8�F2]�J8�����q�������)�oXq��hH�]�9i�eE��x{3�%=c@�LTgY�0ϵ8��2Pʍ�P���*����U��'���N-./=c@�LT2-T��#bYm������*�����D��a�ow��t�+D���l�q���	��>@�h�T&q���g�i�r�rz���xQ��ƛ����!��_K�Yx\��斳���J��^oP�.a7)�r���4GH`�Ώ�o�-nr������k�����~�L���̧th���ħ�l�E�meZݪ+i��,\3DM�`ǌ����m�ebS�f]����Lfg����?*����, S@�����]	M�}����u�>��R��_��H����7uh��F3O�. ���}��Pj���	�`y�=����6�7uh��F3݁��!8�}����u�>��R��_�����d<����֬R1�ɽ�*<e=����*Z�"�#F��8O�^p=���^/a�����6����<���^I=�a-��!�f���v�V8��+ Z����?5�҅7Z���f�}K� �K����6a�s��hp��Ԁ�FjZE��nc�}�I3�-���e���w�\
h�["M6f��������5�JF�M�Vy�cgͼ��UQ�N��V��G���Y���C��&�-�,�X�Ÿ�f�2_B@:P��dS	nT��e�&��F]�J�������	U�֝�%��LP�b�I�hS\'��/���`b]P�L��ϰ�9_��]-͍)�,\���� I���X�%���=��dn'y&̢���N���ꗳ�)�70bxN7~/Ǧ��!Fȵa�E�UJ̘�P���W��-�\��\����WgƘc���Jt���M���bf�\c�ꗳ�)�7�;⑤���a,�"�빱x�Q<�^eg��ɂ����c_�o� x/���C $P��!zsv|MC�[��ĺ6
&���?��������Y���i{\�M�Q#�`>�P����Yy��0�	ĭ��n�W���\?�R�?3�h0)�E�Z��(w
�7`�	�6'�����<5���K�����,%GJ�k���.Ҋ[m]1��F�^v�'-Ɨ�8;�gi��{�]<�S#��B����2"��
��V������+�v��Tj0��L�m��7���dO��H�\?�4x!�i輸m�a��&�^��=3���,je6�����B�g��o&76� ���+ɾJ�Y�WX���v�	p��i���y�6]v��P|Λ#�2�[�k�tf�����0U������J�yP��}H�{_�.�@)1�7-��H�&��_�6�*�q#�L
2�������̹�"�j��;�kԐH`�Q�Cܺ��D�^hא�܇r���+9}�t����{����f�2_B@:P��dS	nT��e�&��F]�J�������	U�֝�%��LP�b�I�hS\'��/���`b]P�L��ϰ�9_��]-͍)�,\���� I���X�%���=��dn'y&̢���N���ꗳ�)�7��y���#H����^'�2����:W�0s�����S�_>gN�-�:'��$+���G(����^Le�0�[��z����jcbb_�B�,��y8f���B6Km���'�5uEq_�<|7.���|N;X�^�I�[\o|�o�����|"ÝW}�utiO����+�%�Q)=d���E@�׺�F�b3��5����4�fgHg)%�RPz
2����$_�>U�V-'�I��.3	
.5�4w���
ק5�C>��M ˶�{T��
�7`�	�6�#'	��m�:��eH��J�	��[W�DC�"�N�?�ot�'��#~D��\��KB����VL��'�s���7K�f*���b�0qK�s��D�1d�	!4wI�o P��z9����D�����e�mu���H��H�
:��p��؋9i��������a:�#�f"�6]v��P��w�	|"�@Ҍp���O��"P)�6�m�`�� P����Y6Z����*y����,��/�&�5K}�*���ՙ��e'�������s�SŠ��z��Qd_No���?�%6=�N����:��*D�)�=��x�Ϟep�h0����p��a!�aG���0������ZT7����:6z��Ӛ�Y�d�.?E�,V z�C�_CeL�f�ZSl�Ȅ�{ڪ0��!�41ҕ�G�9����DC�#�/e�x�P�f��H�H�i�YEK�x7^LX�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�p��vum}}f�|HI�xS��*�=4�Z�P��:M�}���F��E	z�=�Uq+x`\e�ض�,�o��v5ѯ�Ġ�	��� r���] P-I=-$Bf��e�"]mH�ާ��ڣ�qΉ�Ѿ�L��0��p���]y��u����c��oz+�!s�!�9(g�sOwZU��Ŗ9��F�]�����[&u�P\'�L�HoE�AulWD-��V̂�Dw���e�Md^����j�oګZ�Hu���	Ӧ����l�������9)��|{���"z�2�C�a60��P��Ti�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�4)�}Uh����n�r�Z�}=��8��z�S�M:1����oz)���ʠ��6�L�d�[s�	�4�ڟ�Hz�B������B�j�YN")�+��b��i��<�a�]�΋y��%9{��DF��t��-��p�ޕ��M�n}7�{[V������p��ɽ�*<e� ���:H�hy�_��j[�r�����p��ɽ�*<e� ���:��\�j[�r�����p��ɽ�*<e� ���:Ng�2��cD;x�Wp���o�b����RPeA��t1����CԄk�\�!�g�F�s��6���Zr%�����z�:��F#�W��K�_�G]����K�`��
�a��a�a�_��#�|k)&d�BM�P��GrV/Sl�A�B�Z����|�]��w�u��V|`|����2�����jΧ$��Ŗ��'�����䅏�B\0�.�0�	�3A����{'b�T־��Z`�}SG���2�ɗ�D�<䶠�X�������Xƻ�2��D��^��/�����ji�hAU6]?��߇�dG�d��PtD��3;����Hz-yl�:�����Rdst�����j�8]��9r��Z2@���,�o��v./�j�����,�4�����n���8cV�s2����S��-�q��Xv4-��0��N��~����FL��8	�?�b����g�@P�e���k���a;$H{��}7?��yi�Q�f�{��t�����0b��*��-`����g�H��D��[�YA;��<�q�������:�Hb�m{��v].���zR��m�q�G��K�`ږO[})o�ģ�t+��}��Pj�k�\�!�g�xZ�¼�������;A�Y��g����FL��d�BM�P��GrV/S�9�t���P�7ٝGy� �.�Qq�*d��PtD��k�\�!�g��X[�[�*�����Rdst�����j�8]��9r��Z2���-��@L�������[��-�|'Z� ֊�����[,uB,}ŝ�^/aÅ��B\0�.�#�y��T15�T ���ṗ��yw`�}SG��<�q���ّ������?��zF�	D�ܣ{U�荑Z��3������Uj��,Y�^e[��z��I-�C8�RF(Lb����(O%��;!���	��W�Uq f�&�0|5�vUx-��KC�F2]�J8�F2]�J8��� �z F7��2��wz���[g�-��KC�F2]�J8�F2]�J8��o���ٽ�&	u���"�����Ͳ����᥀]a���5����fF2]�J8�$�䠢O)Xv8����9������#�f����И
F�i�ܛ�|�F2]�J8�	C7��3�^��~��Wɽ�*<eɽ�*<e!ՠ��s� b���"������y4�c��)�B=�QpH[��V�H�KV��iI�yl2���ɽ�*<eɽ�*<e�p\�Ì�MlZp
T�m�B���nh��@�;�5����_k`ɽ�*<eɽ�*<e�2+k��˃�6��Rb=LU[$"����N���ɽ�*<eɽ�*<ef3���W��z�2�N�+0C���>MX�1�{��F2]�J8�����q���b�ё�RԱ�-��lb[uO(�П�B
E�=��ʋ5����fF2]�J8�$�䠢O)X�5��M��̠wo�	h�[ɽ�*<eɽ�*<er�~����ac]8���}���W<:K�r�~h8���󞿫�fDq�����yN�F�8I���W<:K#�)L*͌�w�u��V|2�����j΂l�,H_����N���ɽ�*<eɽ�*<eɽ�*<e?@\E��̸B����NI|	*�eF9YH,ɽ�*<eɽ�*<eɽ�*<e�+��%Ɠ�F���]�Ҽ�w	�B�a�h�ɽ�*<eɽ�*<e�����`�k��NL E�២x �ti�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�)V ٥�Dk�z�ʕy��p~rև 낓�q��BE��aꎾ-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)X=c@�LT��q�4Zt6�_� �nx�����=c@�LT��q�4Zt�eif���V�i�E� =c@�LT��q�4Zt`�� �P1s�k��D+;xc&z�j��S�#���%1�M�@`��?�r���SN(1�nr����ˣ�+�������~�1�7 ,D�������E�Zݪ+il�c���k�C �7�W�8+�0�&q���g�i�r�rz���h���*b�e�7�A�&q���g�i�r�rz��[��^Us&L(��hW��l�E�meZݪ+i����n��j�)�5"���R¡�nr����ˣ�+�����#"܇a���[�� b%;xc&z�j��S�#��T6����1QC ��ӑIH���4$�H p~�rj�*���øxQ@Q�;�[U�]Jn��3o�nøxQ@Q�;�,z&�H��=c@�LT��q�4Zt`�� �P1s
����.o`�� �P1shp�|	6��$(�d�z�E�Y0C���>MX�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�YZ͆ˎ����Ֆs?��-��2�e4k|�����in��(����e�c�_?� ���玈��A��kA̍C��4��Ů"�*Q����X���{�>Ə�U�����F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�T�N�:Y�?�ow���I��N�ߤ��Z���`����� NN�d5k2É\"��nr�����].R�{y��z�,U�n[�9����}O�4Ht��Hؓ\\z�E�==c@�LTgY�0ϵ8��)ƙ�7K��)��D]k��ᡵ�	�|pԕzh&q���g�i�r�rz��á*�W��P����оP�E����G�����s�9y�?TZݪ+i8� ���v���x��F���#kN��������C�É\"��nr����˜q�E��@z�,U�n[�9����}O��@��
��)�p��=c@�LTgY�0ϵ8�DfjS��x��)��D]k2�"䊘3��A���&q���g�i�r�rz��(�
W8��G�P���TB�F��w��%~B�W��s�9y�?TZݪ+i� ���CT����x��F�+tT�e��>�U��,��É\"��nr������~֠��z�,U�n[�9����}O��I�%)e��Bl�ȿ�=c@�LTgY�0ϵ8�����+������Ck,�(�[����4j�d�`�"X��S�#��b�Id��}���x��F��!$��փZ0/��É\"������F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�T�N�:Y�?@�>��ձ:����u"��T�
��Z��`��3���x���!rE,
!���"-�o��
���z��@l:s��!�\ `L���,�+���^��w[m�2����@��hY�V�2�ɵ�ZN���ήi�5��Ϥ ��pa�n��Df]?\ڣ�+�� !;�g��'�U�B?|=�Y���^��a�ZQ-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)X=c@�LT�1 ��9���zK�$Ȳ�n�u9{0��%�Zݪ+i�6��#�d];��2ن��K�Ѿ��0�3�1[i��zK�w�d�q�Zݪ+i||�D1��5�w��5�B��؝�T���\\�n�Ѐڼ���h����g+f]t./�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�[6+
ߛ��J�g�d��oz����B��U��Hcɽ�*<eɽ�*<eɽ�*<eɽ�*<eԮ�I��.�`�A��j�����p��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e��h���� *���p�T���\\���|>��N~i��&��nr�����UWѯ���?{�����Y1� ^j�!4���"nr�����lC��f ˯nkB�JMD:�*⹽�H��NPxP�rB	WH��D���ts���K� 0�.{yם�5�^��pj)�0�V-q��S�>¹��r~�����5��I�A���[��Ƹx���]L�E��
����"���M>��USm��]®�,xa��yO$�,�ce���7	��l��6;?;?� ˯nkB�J�,\�le%���u�/���A-�����8�`�A��j���h����]NL��=KT��%z��t�W�\,�5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��� �z F7��O���횑v}��m��ҏR�� f��V3Ǣx�K�-h��($Zm�5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�M-�	zt���u��_a������ɽ�*<e6ė(�t6��Wm*�����Q���X�Y6�Nd"�O���bvz�*�>�������^/a�KW1v�0�2G5�td'QZv�i��`MlZp
T�m�B���Q�w_��T%�3E�|����v��{�����of��Z�91�����<���^ثK*3�Ғ�U��]��`�� �P1s�\�nU^�k�\�!�g�V���P!E��7ۅ���A/��7A� �*C�?�^I3Bv�1��K�`0�G8�rdC��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q���\>ڡO�K|a�� 4��������~��=�� 
��z �W*�D��|F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^��YH1����Ҝ��fat��}����u�9ݓN���˿�ID�b�~�Wr�n �u�HYוۏ�.�E>2�<U,3��ږ����Fnv;�V�
%��
Y\�er"�꺯z^Q,�'�����Q��A��|H�4��b=��K�X�k-­r�wܜ.��dO��@��懡<*h�����1ɾ��ܵ�	5�N���@D�BJ���?�S%����3����V�uCM�1ɾ��rY��ߺ�i�����m�����V�uCM�1ɾ��A �=O5a�����m�����V�uCM�1ɾ��� �!ϑ�cp4`�к`|����2�����j� �Y�\Y�5��y�)�"Uy��\=�B��YX����p��!��E��"]�����;�Y��##A�Y��guDQ�15�T ���`|����2�����j�f��������`�-���Ծ�`�� �P1s�DsF �5�$(�d�����P���H��Q�c���,4���?wX�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�T�N�:Y�?4��!��Yo����d���^�͎��VJUT���K��
6ҹ������c�D6 �z�2�C�a6
X��`��~�b�b�	�� !;�g��׊KW��*�D��|F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�0C���>M����sv�k�D<�P,��D�����a.E�O��ʈ�T+�)J1�tM�|@�ĩi�]�C�F$�aD��4>Pܓ�O���PGkPl�ޛfe�^C�ɽ�*<e[�Q,�o��v��c��/eJR�k�!�����,ɽ�*<e}��&�rSV7�@3�w�K�Yc��� Nb '��D�Lg ��ۘ�(��o��_o��u��<_��iM��=~"@��[f/������$�6g��xy� Z���7�Pa}��I`��x"��W=��M�,�r
��_���׹��wl��k���,(nɽ�*<e2�����j�-�On+#�M�mZ ������"Mɽ�*<e[�Qpx��������H
��oC���SMWK5�ޭ {�LGP�P�7ٝGy�YZ͆ˎ��_�bOh���5�T̬ϭ�D�����a.E�O��ʈ�T+�1w�s"���_�J��]�C�F$�Xbf'�����Ҝ���	j�֏�x{�������p�������`���K�`�V�G�j�U{]%�K�P��mɽ�*<e!��E�q������'-hpG����p�q^�/�D���8�!�|9�ݞR��=�˙w�:�G14$���)AU��v�r@~h�,�{m�:V��~���:�7���?�K��wx#T|���*!F�B�� {;�3-�Q-K0qt�E�x���]L�Eɽ�*<e-��E)�VAD���9&�v�J3�tMB�]��������p�������`�-���Ծ�`�� �P1s�DsF �5�$(�dؤN\=�P�7ٝGy�YZ͆ˎ�}*��2�UްBL�f�XY��D�����a.E�O��ʈ�T+��BW�2@�	�x��`��]�C�F$����r�r����Ҝ���	j�֏�x{�������p�������`���K�`�V�G�j"M�VyQ�K�P��mɽ�*<e!��E�q������'-hpG����p�q^�/�D���aK��N9�ݞR��=�˙w�:�G\?��;(�G�8(�6��r@~h�,�{m�:V���G�A4P�(Cԑ�r��wx#T����FcZ�B�� {;�3-�Q-K0qt�E�x���]L�Eɽ�*<e-��E)�VAD���9&�v�J3�tMq>{�f�/����p�������`�-���Ծ�`�� �P1s�DsF �5�$(�d�����P�7ٝGy�YZ͆ˎ�u��NEk#Z��v�ŭ�D�����a.E�O��ʈ�T+�ZX��f��Nk�z�9�]�C�F$����</�m2����Ҝ���	j�֏�x{�������p�������`���K�`�V�G�j1y��1wjVK�P��mɽ�*<e!��E�q������'-hpG����p�q^�/�D�6��n9�ݞR��=�˙w�:�G����w(c�̨T��N�r@~h�,�{m�:V��tXƐ�p1���#���z��wx#T8�r���B�� {;�3-�Q-K0qt�E�x���]L�Eɽ�*<e-��E)�VAD���9&���fݱ ���(�r������p�������`�-���Ծ�`�� �P1s�DsF �5�$(�dat��Y-��P�7ٝGy�YZ͆ˎ�D}DQ�*q�H���A��D�����a.E�O��ʈ�T+��ܢ�o���F�4����]�C�F$��e< g�\����Ҝ���	j�֏�x{�������p�������`���K�`�V�G�j��I�,�Z@K�P��mɽ�*<e!��E�q������'-hpG����p�q^�/�Dm�̓�D�)9�ݞR��=�˙w�:�G�ڒP%��%>Ʈ��r@~h�,�{m�:V��jK��z�_a�L��N]��wx#T�	����B�� {;�3-�Q-K0qt�E�x���]L�Eɽ�*<e-��E)�VAD���9&�����ḵ�(�r������p�������`�-���Ծ�`�� �P1s�DsF �5�$(�d���K�KP�7ٝGy�YZ͆ˎ�ҥ�53���M �r��D�����a.E�O��ʈ�T+�b��lL�ic�t����eN�\"��S���`���`V�f�Bɽ�*<eV�D�=~�@L������U^��#��U{]%��NSad���p\�Ì�47��ט�@��p�q�nvo��c`�� �P1s�lT�P����_0(I4�������*�R7���ΫU���0B;�㶛�Ĉu�"��1��IS��}.3!LZ�Ug�7SM��wx#T�����d�x{�������p�������`���K�`�[�Ot=�;/eJR�k�K�P��mɽ�*<e!��E�q������'-hpG����p�q^�/�D��+?{B�JAj����x �J8���5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^�����j�Ԩ[��d�V��{|r[�i']n�u�U�i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q������2�f3�I�^S*���������ظ5��Oh`ò��O�e��^#G����p��� �<%@u�\�1��/nɽ�*<eJПE�[5ɽ�*<e��ٛ�ɣ�����p���_����i(9RV��9�pɽ�*<e[!]��{H�TωnJПE�[5ɽ�*<e��.t���90��Z[����x��F�Y>u���kɽ�*<e����@��G�n��0C
�V[�'$��R��e�����kV�f�{��t���FLE+����kp�l}Rk!�|F͇�*�����r��s(�?A�Ҏ&�Ё?m�-�,�X�Ÿ�f�2_B@�~%.DI���:��t�%2�/	J��hא�܇*9�2�\c�5��u|R���GX��a��Xڟ3�8�H�d�h���� I���}�t�wI'[]
*�J���oE����:��C�$k5p!,�7ڐ9� ��h��'i沃�Z}����Hc�9�%�\T|Aů� �B�#��t�(a�����z}�E!Ͽ���!Lؒ&�bL�.��. ����lB��,zyj���0_��A�\��B�N��%졖*��j)?��(a�����@��$�G#�ӵI�0��#Ҟ�s�-I@>������BP�\_�0'���I"ʈ�W�rB�������i0aXK��2��H����D���i�6 ��Z�)a��\ `L���c��}W�R�#C,��n�Yx���|��/_��P��r�k���g��� H]K�s��K���{T��
�7`�	�6�#'	��m�:��eH��J�	��[W�DC�"�N�?�ot�'��#~D��\��KB����VL��'�s���7K�f*���b�0qK�s��D�1d�	!4wI�o P��z9����D�����e�mu���H��H�
:��p��؋9i�^��,1DԾ����\J���H�.'a:�s�c�A �Ы���VI#�1z���x�q��Ǝ�b\[��½�#��$̆���5��0^v�'-�r�D��6�^i~��b!�t�&��9W����m�$��mtM#�/���g���x �&�����GX��a��Xڟ3�8�H�d�h���� I���}�t�wI'[]
*�J���oE����:��C�$k5p!,�7ڐ9� ��h��'i沃�Z}����Hc�9�%�\T|Aů� �B�#��t�(a�������bc+Ji �8s����6e���%���2"��
��4N;L�Oc]����m���x�?���wIF��E��OU���2ޔ��e�����{�n�q�r/<��\�D?('h(�m�W�K.j\�NIf���'Q+j���p�D;&��'��K�����c�׈�}���	'��@Ybs����Q��� ��ɬw��2,mD9���\��w�0��8w���c�Y�l�%�tB�;��Ha�L�zַ��-ro��S�7>�<S@��9jj ����̜�ߑk���g���>�0 ;��od<~R��Ǥ����e�9�\?%&�/�~=rN��uL�7d̈w�U���YEL8��L�Y���ay\�n ���J?|��'�[����K���3��h�A5�oD����S�_>gN0e�,F��Т�����[���ɛJ�z6Ǡ$^�H�#��]G� ��\J���H�����v\�k�tf�����0U������J�yP��}H�{_�.�@)1�7-��H�&��_�6�*�q#�L
2�������̹�"�j��;�kԐH`�Q��
I�DYZ�?�0.܍�G.I�TVzi C�"4D�MUP\�0W�1�5<�蔺Z�ØKϿˬ����B�Vh��lk�D�`�wQEE�,ߨ0�iN�x�*B��0�ѡlv���tk���I���v�D�t*�gc�꺉�@jB��Z�!�W�/�Cd�سy�%�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S�?%6g?��U�ӕ'�j~��fvF|RD����nfE]�l�VH����-ʀ?� 8�\�/k�����P��'<�",
!������W824��o�v��� !;�g���RH��.�"��.�1�5��P���p:��O$b�����9.��7Ļ1"�p<Z���X$���L4�DكV%{�v�7��������7�����'��R�@	�#�i�z�~@^T�'VR ME�99^qy�t�(Y��ex�j'���v�ϧ13��K���ǋ_��k�� Ge�[��T�˚�j�X�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��"�iS{/E�́7�׈�|�.�Q>���ě��Fnv;�V�
%��
Y\�er"�꺯z^Q,�'��ƭ26���\�����R��dL:����2�����Q�k��/�� ���:Y��$C(E�Hw^���ɽ�*<e�TwR��U�{������1�ˉhύ.P�ɽ�*<e�TwR��	bV׶X�׾��1�ˉhύ.P�ɽ�*<e�TwR�����d�on�[;�8߰+,���h�!��q�<䶠�X�� �*C�?�P���H��@�D۬�}~�a�h�!��qM�
��.m���Y��؛rY��ߺ�iA�h���f����N����M��L׆"�@��D)�#�y��T���`.}���W<:K���K�Js����t�~G�@����ƚ��U�H���jp����FL��[�3���z�2�C�a6i����hB��L�f�y}��Qe��P$4k�DQ��t1����C�qbaZ�4Ow��g�.Sk�&!6�]{��}7?^(b��n9%���vc[���%#�`|����mv�Bӝ`Z���#dJ)N���T������Q�`|����2�����j������;��_0( �L���y��W8 �+N���ط@���z���J)�����K����7���^/aÅ��B\0�.U����,@L�������[��-�|'Z��hAU6]?�2�\���2pG�Z?)���g�H�1j��2��C0M`�ܙ)w撨�fx�k�dPY��$C(E�&#��y#\�5!��s�*�V���~f��(`�Mʥ����w�'T(��Î�HX��`�+t��P���.,h,�o��v./�j���^/aÅ��B\0�.�#�y��T15�T ������L���1��0���g�q\��#�H_�s��0�T[�mv�Bӝ`Z���#dJ)N���T������Q�`|������<�K��e���k���a;$Hb��������)D���A�Y��g����FL��d�BM�P��GrV/S�R�c�Mt��&
qy��fx�k�dP#L��0����ɖY׎�+W���%#Y���L}Rk!�a�����~�݈����;�r�����׀t���8ο�K�����j#�HS�� EYZ͆ˎ�F2]�J8�F2]�J8�T�N�:Y�?XF�P��V���/��YZ͆ˎ�F2]�J8�F2]�J8�T�N�:Y�?J�ۇ�5�!o��c��Q�-I��a��.�+:-nP�����F2]�J8�~�&T�S��)`�"����
��䭍����3��B
E�=��ʋ5����fF2]�J8�$�䠢O)X�yl2���ɽ�*<eɽ�*<e�p\�Ì�'�09k� ����>��y~��P�  �g�l�O6d)8�����#��g�^5��Oh`�wo�	h�[ɽ�*<eɽ�*<ec�XO�_ag�̸B����NI|	*\�I;���ɽ�*<eɽ�*<epH[��V��"vЅ\�P�TT�I���W<:Kɽ�*<eɽ�*<e!ՠ��s������V<�κ��_i�ܛ�|�F2]�J8�	C7��3�^20p{>}.^9j/���B�4��,��s� "m�r������F2]�J8�~�&T�S�ic��ݤ��B�a�h�ɽ�*<eɽ�*<e[�Q�=��c��v�5��M����Հ��-Nc'�T?�������VL�H�KV��iI�5��M����Հ��-Ncź9�/��-��E)�VAA�h���f���W<:Kɽ�*<eɽ�*<eɽ�*<e[�aʎl���!�(I�=LU[$"����N���ɽ�*<eɽ�*<eɽ�*<eщ�N�#�9V8��+ Z�"�����.�^<�
:�ɽ�*<eɽ�*<e�K,V[dM'6/�`�+����5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��� �z F7H�(�O(qb�R#l�Bq*�{{e���5bYZ͆ˎ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S��H p~�rj�*���øxQ@Q�;�du|K�H p~�rj�*���øxQ@Q�;�~��5!�H p~�rj�*���� Nb '����@WW���������Zݪ+i�sk�=�ߟ�@� � �e����x\��斳�w_��V�J�k2���z���ob!,�1v�w�ow���v��}�]=S�Z�:��C��>M��;xc&z�j��S�#����8xyb3�lK�,`�;xc&z�j��S�#������S���hs��#f5Ҫ���ow��H���?Z"��f��(����/=��x\��斳�w_��V涾����� �缬��Vu9{0��%�Zݪ+i��,\3DM�.�E>2�<UR��Az��&q���g�i�r�rz���USm��]�g�Xy�6�«&n�U�USm��]¨��ҮE�H p~�rj�*���� Nb '�Φp�\��� Nb '�k#���IY����H
�ը��ҮE�>&��l-�i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�)V ٥�Dk+�&�<�C�
�jӁٗL�ߨ����^�i�K��=�%��!�/�'fh�hN�����F`F��� �=H�|��G��]�S�[��H��=�b�C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q�݊����F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�T�N�:Y�?@�>��ձ:����u"��T�
��Z��`��3���x���!rE,
!���"-�o��
���z��@l:s��!�\ `L���,�+���^��w[m�2����@��hY�V�2�ɵ�ZN���ήi�5��Ϥ ��pa�n��Df]?\ڣ�+�� !;�g��'�U�B?|=�Y���^��a�ZQ-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)X=c@�LT�1 ��9���zK�&�IòG�;xc&z�j��S�#��{�����Y1� ^j�!��s�~D>K�c�5������m�;xc&z�j��S�#���H��NPxP�rB	WH��ߖ�on�������)���k%J�?�USm��]�݀F_zT�ɽ�*<eɽ�*<eɽ�*<eɽ�*<em�!Z2�e];��2ن��Z��V�O����ɽ�*<eɽ�*<eɽ�*<eɽ�*<e���<�&f�:~�)=R�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eɽ�*<e�USm��]��,�t�l~������)u�g**��],����ow���;�
(lx�@���L���9�<Ѻ�;xc&z�j��S�#��%�y]�v��G��̿5���caګ��8�����|��h�����:'�L�7��(��m�� Nb '��P���;݌*�`Փ��[��L�)�����F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�T�N�:Y�?��5	oU++P�]�q���U�H����3SY������S����8{�F������F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�T�N�:Y�?Gi
��Cj��I>/�4	(yaf��ٿ	�����qn�\DԷ��J}��Pj.���8�j�<�U�q;��N+ށ��P��7M�}����u��Y�#�&�����d<�2�>��1c�XO�_ag�̸B���ثK*3�ҒGi
��Cj��W���#��U��Z����˃�6��Rb�����E+��I�ź9�/�闄k�\�!�gi�.�!/��o������/��K�k�I9^�ï�Lz�����K�P ��謋:��5���ڵr�����(RZ^�%?J��,^��%�[�3���Hf��1��Gy6+�$��ٜ�N�� Ge�[��T�$�)o76�끆E�n`|������<�K��H���Ck�끆E�n`|����jy��0Dφ�H���Ck�끆E�n`|����2�����j�R"'lvsJ�>�z�{���[���MĞ�1�ys���qk�N*�%�Ir=Xl���`V�f�B�p\�Ì������7;��N+ށO ��sye�ɽ�*<e2�����j�5�4����>�z�{���[���MĞ��c�R��-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��l��q���S�l2��@�D�3��7ZK�[��M3)�$N5G �):B�RtnGP��'<�",
!����^�I4�(V>9��DkQ6�Qod|-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��l��q��&5�_�vr���4GH�n �u�HYq�����0ilw|����Ω��Ez`r���AYmu�O�
�����+x��o��mq�͝*�x���]L�Eɽ�*<e-��E)�VAD���9&���C�Օu:׈S�yß�Q{u\�0C���>MX�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�T�N�:Y�?��-��'��[�y���ۓyP��YZ͆ˎ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�?��F�-��C>��M �IꜦ��/�����eA�Y��g��~��W[�3cX���!D��'�vS+ё@n1���Or�/~r�&V\
���|H�Pk���,(nɽ�*<e��u�<6�ɽ�*<eK�����h����N�ߔG�=��r��W�*�`ϭrV7��<_k�k���,(nɽ�*<e?��=��5�9���S\_@}���^��gƇ�e�ɽ�*<e�����I��rc嫨��~����p����8t������p���+�r��y�=����lQ+�or��1��������{9���i�O��n�:Y�f�H3UU���f�O@g�IFS�w�s@�����4�
�����%nġCB�I�t�`H�Q����U�xl�(T�W#�(�*� �.6p@�*3d�#_�0!s�,�	���
6�.8�0�T��(�H���-)�|�d!d�H�d�h�ݔ�x��{��õv�̟��������.s����g ��$�L��ow(7ALۗ)��/��	`�)�h��{̠����Lʉ/[¶���`���c��� �	[�w:���ע��������t��E�̎����D�<L}ڈ�����dn'y&���3��ͨL���K��a9q;���]��e�G<���ߤ#����ө�((|�w��M{� C<�ls���|����䋇�æ��tg������a��4W}����Y[A`�_Z_MyV<tn�||oKװE��"
8��o���l��͡U�R�4�t���#,�>�Y����,�:�+[��epՈI��	n��WO�.�<8��]���f8��H�\J����K=҉7�#������g~�nR�&x��l���Hwa_i��\{��ЍM�Cʌ���H�v���5������A��\��G������Oc]����s��� �F��.�8X��)8�\/,AܥЍ�ө�	I�\���YVeX���V�E{�49��������4�=z��F		DAu��6YhzoC-x�i���
V�r&A�V�6�.j���|R��Ǥ_�|�P��L���Xj��)�*��e/6�5��0�K(8 �%D\������A���UJ�l�t�p,|4�^,e�I��ހVh��rd�#�®c��P]c_��g�k
�G���0��'����u����<LO��$����tk���}Ո�,�AQ]�h�j�v���� ��B迅9DԄ�r7uo)V�&�>\���^��0*eL���J:Գ�5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�p��vum��^�.h�%Ѷ���\��fvF|R*o��A���^�2W��@��:M�}���F��E	z �2B��"KD��%�+���9 
HpT�t��E ���L7bZ?����@&F2]�J8�F2]�J8�F2]�J8�F2]�J8���ա8&�o�	rr���6�XoN�L����A�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8����b�bgxP�8Y�R#l���/���?�pأ�a\8�,��/�p+�3���^������eX�3%7|P�̖F��xg�t�2M�b��i��<�a�]�������P{���R�B��ɽ�*<e�c;��},n�*��g�����8�ɽ�*<e`�w�A���?���3�
���=H��Q736k�:�s	Kz
��NXWɽ�*<e������o�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�S<��1���F2]�J8�F2]�J8�F2]�J8�F2]�J8��<�2��M%mD*��+�G�O��d��[�u�aH��[�ї'�h02%Qk!F5ğ��ه�rݶU���e�y0ѷ��h���9kZ���v�t!cJ(�Z�0�W4iE�a�Q�e:���,�	z��$�P~F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8����Ѹ��:����oz)���ʠ��6�L�d�[s�	�4�ڟ�Pc.��P� J�F�{��8B`}���^b�AaKC��ଡ଼�F2]�J8�F2]�J8�YZ͆ˎ�0�`��D�����F2]�J8�~�&T�S�5��Oh`��B�3�a�6��mL���$��J� ���	/5��Oh`��a�u R���^7��L���$��J�ԾbQ�����ºU����6�/G���5��Oh`M�p�+0�{��:��$B9Hl�+s�z�g�-L�����S�4(8��pM]�Ҽ�w	�B�a�h�ɽ�*<eɽ�*<e�2+k�ݠ����d<�s��7Z�yl2���ɽ�*<eɽ�*<eɽ�*<e��,#D7��K�am@��r�Zjsp�6?���:�ɽ�*<eɽ�*<ef3���W��z�2�N�+0C���>MX�1�{��F2]�J8�����q��U���'��|�~���Ǌ����F2]�J8�~�&T�S�ic��ݤ�����a3mɽ�*<eɽ�*<ev�L{Ǘ%>� ���	/ic��ݤ����l�*����}I����nX���ʚ���&
���b���$7O����h���?K����9�֣��K�Js���a����+��K�`� KЋ��>R}9��V+#�yb�����N���6����=�ɽ�*<eɽ�*<e�������!�(I�=LU[$"����N���6����=�ɽ�*<eɽ�*<e��$S�(���K�am@�nh��@�;�5����_k`ɽ�*<eɽ�*<e�p\�Ì�旿�]���6�z�������F2]�J8�~�&T�S��)`�"����D2x]��S��pľ�ߊ����F2]�J8�~�&T�S��x���z�k<'����	�����?r
�x�1;����yf4�H�+_8�,���3�d=�� �;�"�<�*ʣ�Pwf����XS����[�A5��Oh`0ZI����L%V�
������/b�r�m0{���N>�j[�4�U.�
=�������)�h�s����K��e=3s#�/�;fD�/�Y��E�Ի��(f�@�~�K]�Ҽ�w	�x�Ae�+S�Ξ�����x\��斳��Y���fK����[1�W_K�Y��{v�����?���3�<�&���t�6�Z�З�o\ע����g��5����fF2]�J8�$�䠢O)X�����)0��\���4��5����fF2]�J8�$�䠢O)Xj`▘9��e�=�@侮/�žC������7�!I�2r���4GH�n �u�HY͌r����������7�����d<�2�>��1c�XO�_ag�̸B���ثK*3�Ғv�L{Ǘ%>�"vЅ\��Y�5�8��,#D7��K�am@�p���b�!׈�����7,�o��vr���4GHB9Hl�+s��s�Gv�<���?���3�����t7��K,V[djME���:ɽ�*<e�����g#!x%q��~�U�c�� b���.��ݞ�Z�_o��u��5����fF2]�J8�$�䠢O)Xn����K�pg���fr27�?����i�ܛ�|�F2]�J8�	C7��3�^}��Pj]��w��\��)���� �A�����Y��^/a�zpt�d$\�5���D�8gg:�lx�f8�i�`�1�c��Xv�e���S~Ti�ii�Ӄd7۠+)�Ay]��rO����xŗBGj{=E��Rxt��(�^X��yO]�&��I���R��A|`�$������kȡ�B,ŭ_
j�����ͬT$OeMS���s�C�罤�9.�f�i����
D��H7����{�ƥUuh��V�g5D�l��9q�X�:׮�5:��KL����z�>�4[���{u�^ק��}�{�ʘ��SD!��Ю���0�V�٦�����2���X�����wD`֡��y����"�m���F^��`���#H����^'�2����:W�0s�����S�_>gN�-�:'��$+���G(����^Le�0�[��z����jcbb_�B�,��y8f���B6Km���'�5uEq_�<|7.���|N;X�^�I�[\o|�o�����|"ÝW}�utiO����+�%�Q)=d���E,��h��DZ�x���F\��w�0��8w���c�Y�l�%�tB�*��� �&&s�:v3�9?k����Q������L�����p�N_�qe�
��>̊��%�
�T���k���g���*�F/��q+�\��$|?G��a�G�x�D�9ϑm�eQ���9*Q����� P�7+��$-���G[�z�A��ie�\#�_Hc����'d����uC)�E���Q�0)Dm*
kma��ݑ�`��N��X5/�)I�|��o9�H[��UF�n]h�^�o��p����=����+P
���(�5;B�W��M��v��E�`�w$�P��j�:�mheˣ��:��?Dg,2ms����{Ue#T&�ީ�q�� B�����z"3�������kȡ�B,ŭ_
j�����ͬT$OeMS���s�C�罤�9聯�v!�������k{��Ty}�zj�"��0��U��j )���.s���2D��%_�y��N�[\��NT��>n.r�P�S��И]h����,��D�se��L���Ӡ��B:l��9q؟��?��6\F�߉�}3z�s"�!6���f����!Lؒ&�bL�.��. ����lB��,zyj���0_��A�\��B�N��%졖*��j)?��(a�����@��$�G#�ӵI�0��#Ҟ�s�-I@>������BP�\_�0'���I"ʈ�W�rB�������i0aXK��2��H����D���i�6 ��Z�)a��\ `L����B)JǴ��	ĭ��n�W���\?�R�?3�h0)�E�Z��(w
�7`�	�6�����C��F���Y��U��>��M���2�أ���Q������L�����p�N_�qe�
��>̊��%�
�T���k���g���*�F/��q+�\��$|?G��a�G�x�D�9ϑm�eQ���9*Q����� P�7+��$-���G[�z�A��ie�\#�_Hc����'d����uC)�E���Q�0)Dm*
kma���t�jp�]$u�	8'��v�eMV�z�U܉����4�=z��F		DAu��6YhzoC-x�i���
V�r&A�V�6�.j���|R��Ǥ_�|�P��L���Xj��)�*��e/6�5��0�K(8 �%D\������A���UJ�l�t�p,|4�^,e�I��ހVh�.v�#?kS�x���{��I7�������j){c��P]c�1�\�r; ���ڶ�du��όT(ɇ�qkaDt¨���:!�6AD6B�iٲc�z��+��+T��L��l�����O�l�[#�e�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�dPؔ�(�{ԅӽwA�?ӡ�M�ጋ5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�
�c���z��g:�Bح������A�Iԗ.*�ȋ5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�]^�h��/Uz	��� �'I�F�IGzB�r�J��9WQ��,D������8��7����ʠ��6�L�d�[s�	�4�ڟ�BZ;�(}�}�O�ɧ���Ɯ�hy[�6p��WS�X��"�W̌at�)�����d���l�/zɪ�퍑I�a����̶��&p�����&p�����&p����@<��l�be�a�i|������PA� ���NHI��5da�Y)(�[���3��/s!_ǁ�y ����IuW��;+�%��$�]}0كG=ͷ�@�������W��Ԁ��/��<�����L�w�h���*b�:��Jx�C4�#�y���|��m-���)D����ά��������KxX�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�^��'[�EEѤD����8�3�F�K2f]}v���^B%B����ŋ���l���8B`}���^b�AaKC��ଡ଼�F2]�J8�F2]�J8�T�N�:Y�?2����>YZ͆ˎ�F2]�J8�F2]�J8�$�䠢O)X�yl2���ɽ�*<eɽ�*<e�p\�Ì�D�H`4�!G���R������x�17�=p�J�滋��׿o$��^�]�Ҽ�w	�z�:��F#��\�{[��5� 2�9�l�,H_��� ��#*ɽ�*<eɽ�*<ef3���W����BV��xV8��+ Z�"�����.�^<�
:�ɽ�*<eɽ�*<e7uh��F3˃�6��Rb=LU[$"����N���ɽ�*<eɽ�*<ef3���W����f�}Kk�y����5����_k`ɽ�*<eɽ�*<e��0�(��� ���	/5��Oh`)���Q����v��x�\��b/]�g+:ȅ�J�_���G�P�!R����R�nhs;J6'���]�Ҽ�w	�B�a�h�ɽ�*<eɽ�*<e1|g��2�>G5�td'P�TT�I��~��Wɽ�*<eɽ�*<e!ՠ��sd+r9�N�Փ�F���M��1����.�^<�
:�ɽ�*<eɽ�*<e� ���s^q&/h.�yl2���ɽ�*<eɽ�*<e�p\�Ì����=�D��G���R������x�17�=p�J�滋�ƨ��j���]�Ҽ�w	�z�:��F#��\�{[��ԃ.�n�l�,H_��� ��#*ɽ�*<eɽ�*<ef3���W��%�Qx��V8��+ Z�"�����.�^<�
:�ɽ�*<eɽ�*<e1�o�5+�˃�6��Rb=LU[$"����N���ɽ�*<eɽ�*<ef3���W��<:��y,4k�y����5����_k`ɽ�*<eɽ�*<e���� C��� ���	/5��Oh`)���Q����v��x�\��	�ݣ`ȅ�J�_���G�P�!R����R똁F"��d'���]�Ҽ�w	�B�a�h�ɽ�*<eɽ�*<e.d���d�G5�td'P�TT�I��~��Wɽ�*<eɽ�*<e!ՠ��s�A	��r��F���M��1����.�^<�
:�ɽ�*<eɽ�*<e=/�lx�
s^q&/h.�yl2���ɽ�*<eɽ�*<e�p\�Ì�ڂI�j�mG���R������x�17�=p�J�滋�ƀJ�k���]�Ҽ�w	�z�:��F#��\�{[�z��/Kx��l�,H_��� ��#*ɽ�*<eɽ�*<ef3���W��;�W���<V8��+ Z�"�����.�^<�
:�ɽ�*<eɽ�*<e�Z�E�I˃�6��Rb=LU[$"����N���ɽ�*<eɽ�*<ef3���W����z.���k�y����5����_k`ɽ�*<eɽ�*<e����h�+l� ���	/5��Oh`)���Q����v��x�\��ϰu��ȅ�J�_���G�P�!R����R��y�H�6�'���]�Ҽ�w	�B�a�h�ɽ�*<eɽ�*<e��&0Z�G5�td'P�TT�I��~��Wɽ�*<eɽ�*<e!ՠ��s�RE��и��F���M��1����.�^<�
:�ɽ�*<eɽ�*<e�����s^q&/h.�yl2���ɽ�*<eɽ�*<e�p\�Ì��C���<mG���R������x�17�=p�J�滋��&_�Z]�Ҽ�w	�z�:��F#��\�{[�	rU�O�Ȃl�,H_��� ��#*ɽ�*<eɽ�*<ef3���W��Ǭ�U�V8��+ Z�"�����.�^<�
:�ɽ�*<eɽ�*<e$�F��˃�6��Rb=LU[$"����N���ɽ�*<eɽ�*<ef3���W��v�Cr
?�k�y����5����_k`ɽ�*<eɽ�*<e�T;�m�� ���	/5��Oh`)���Q����v��x�\����ȅ�J�_���G�P�!R����R�[��mB='���]�Ҽ�w	�B�a�h�ɽ�*<eɽ�*<e����eg(UG5�td'P�TT�I��~��Wɽ�*<eɽ�*<e!ՠ��s�X�k�9.���F���M��1����.�^<�
:�ɽ�*<eɽ�*<e	�=�fqs^q&/h.�yl2���ɽ�*<eɽ�*<e�p\�Ì�_�@�w��@G���R������x�17�=p�J�滋��_1�|y�8]�Ҽ�w	�z�:��F#��\�{[��+�������l�,H_��� ��#*ɽ�*<eɽ�*<ef3���W��[Eu�3/@V8��+ Z�"�����.�^<�
:�ɽ�*<eɽ�*<ed��8�X˃�6��Rb=LU[$"����N���ɽ�*<eɽ�*<ef3���W���x�Gᑻk�y����5����_k`ɽ�*<eɽ�*<ef�{�먕 ���	/5��Oh`)���Q����v��x�\�\�j�l�ȅ�J�_���G�P�!R����R�=|���w'���]�Ҽ�w	�B�a�h�ɽ�*<eɽ�*<e�&k'�|G5�td'P�TT�I��~��Wɽ�*<eɽ�*<e!ՠ��s���+��P��F���M��1����.�^<�
:�ɽ�*<eɽ�*<e9���&���s^q&/h.�yl2���ɽ�*<eɽ�*<e�p\�Ì�P���U8����k�L���G�P�!���}I���\�{[����O�U�u�(`h���8���.�/)h��Y#�ؑ�b> |�!N5��Oh`�wo�	h�[ɽ�*<eɽ�*<ev���[eG5�td'P�TT�I��~��Wɽ�*<eɽ�*<e!ՠ��s����@a�V8��+ Z؋$��,!i�q�k�אɽ�*<eɽ�*<e���la@:x����Q��]�Ҽ�w	�B�a�h�ɽ�*<eɽ�*<e���-e��=��c��v�yl2���CCgm�0�w}���H��=(�%�ʥȅ�J�_���G�P�!R����R�2�����K�`�"�����.�^<�
:�ɽ�*<eɽ�*<e2���"�#F��87U*���g5��Oh`�wo�	h�[ɽ�*<eɽ�*<eJ�H���N���<���^�NI|	*�eF9YH,ɽ�*<eɽ�*<epH[��V�vt8�@�J��;-��+~�5����fF2]�J8�F2]�J8�)V ٥�Dk��dń/0-��KC�F2]�J8�F2]�J8�	C7��3�^���W<:Kɽ�*<eɽ�*<e�K,V[d[g�R�mM��1���ۏok|� �|�T+���-F�s>-ʾȅ�J�_�����N����M��L׆"�w�� ��b> |�!Nic��ݤ��B�a�h�ɽ�*<eɽ�*<eȌ���\�m�B����r�Zjsp�6?���:�ɽ�*<eɽ�*<e�-���*����<���^�NI|	*\�I;���ɽ�*<eɽ�*<e[�Q����6��9-��KC�F2]�J8�F2]�J8�	C7��3�^��ՈW)��MI:��+�BuK#[i�ܛ�|�F2]�J8�F2]�J8�]�Ҽ�w	��f�jd�p5��Oh`B�2>��w�d�q�Zݪ+i�?�7��5S˝�#F4��qլ�17ӹ�qDy��l�E�meZݪ+iZk���"�#L-�qo�7y�i�t�1&q���g�i�r�rz��v�Hn/��Be�5E�k_K�Yx\��斳G��_]��Y�!9@�73q��)�U@mu9{0��%�Zݪ+ix�[H��6{��tr�Ɉ�qլ�1;xc&z�j��S�#������S����n�0���#Wa���H p~�rj�*���\�`�P�J��wP��9�ی���m*�D��|F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�YZ͆ˎ�3VU=f�:>-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�_���9�fYo�u�0��zl#�D�>֠�E).��О���}�;�ߠ�{v���.4%�X��҇�s�����Y��`d��\�Z��?�Vl��nj��K���{n�AW��A��:��$�ur��!�N�
�I���o�u�0��zl#�D�>֠س�H����T�Ê
!���2I��j��K���{n�AW��A��:��$VG�X�y�k�8@��z���2I���)��Q�Ϭ�'�5��{b��D�[�Q�_x�'��E��7ۅ��&ꬶ�Rɽ�*<eɽ�*<e
1����+�6�I�]'E���iɽ�*<eɽ�*<eɽ�*<e6����X�(*�
�x����gI�N�ʆQ'�ɽ�*<eɽ�*<eɽ�*<ep�t�ƍB6G4���E��7ۅ��b�-:�x�Q��>�zf� ������Y�ǭ:9���Z�!��2���C�sNq�0a�E�I�����}��_x�'��E��7ۅ��b�-:�x�Q��>�zf� �����쓪?�� ���Z�!��2���C�sNq�0a�E�I����:%����ܗ�_x�'��E��7ۅ��b�-:�x�Q��>�zf� �������0��݊.��Z�!��2���C�sNq�0a�E�I���䞨��)���_x�'��E��7ۅ��b�-:�x�Q��>�zf� ������%�{���g��Z�!��2���C�sNq�0a�E�I����,�2���_x�'��E��7ۅ��b�-:�x�Q��>�zf� ������<o/��?,��Z�!��2���C�sNq�0a�E�I����z��X^�Y7�_x�'��E��7ۅ��b�-:�x�Q��>�zf� ������\O�{�؋74����ɠ�{v���EQ���ߓ�,����nJw�s[zc��Q�u�w��"��m�
9g�}�zLW��~��j�B����/E��+�(�T	��(�[�v��ǭ1Z]�/���JH�I�6S�@��#2����?5���rݯ�����B�����>-���<�WV
v������Q�}ؿś��4�;����>�������^/a��]�p�p�f��.[��N��[QjJ�L������a�+R)$��Ι��BAw�R��;��2��:7}��Pj��^-4�&%���u�/�67�lȿ�}����uoҲ�j�U܉��ܫͰt�H:�4�1RMQ¥�g�}�zLW�:,���ϼ)�KU#i�+�(�T	��(�[�v��ǭ1Z]�/������ۧ�}>�������?5���rݯ��tĕ5�!)k0�[�+�(�T	��(�[�v��ǭ1Z]�/�������O9)N��5��S����?C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S�-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�)V ٥�Dk�%a���n# �
����y*�D��|F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�YZ͆ˎ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��O��e��q�\z� ���zl#�D�>֠��~�;5��'4M���/v`S^!����������/TB����/E�6v2���A�Y��gį�Y|����ȁ�\�6v2���A�Y��g!mCd7$w�*j����6v2���A�Y��g���Q�fӔ)L�f�	6v2���A�Y��g�>�u+��;{kI�6v2���A�Y��gğ��Ժ�ېր*�6v2���A�Y��g-�E�L���	�˶6v2���A�Y��g�wF"Q�X'�/�JA�a6v2���A�Y��g�j�{�T�)�KU#i6v2���A�Y��gr��-j;o�diF�6v2���A�Y��g�OA��(NKQ�A��I���~*�Ջ���:W��^�{$��JH�I��ha]���~��7����
�9�����(�[�v��HvК��O�9?<076��~-y7:W���ڬ����_d8��W���{�j���+��m�ej4Mo��}g������+C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S�!�nUrW��/І��4�qC�S��"|�J����0}'A� �����>z�^�9�!���"�O�c������S�y|5h��Ϊ����Gph�����)vX�-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8����4T!��]0;�G�	�M��)�atBҷ��c A�[f�矑��ӆ�澮/�žC���U�8�sl�Z)^��_������w��4�.9���ՠ���l$���I�\!����P�7ٝGy��ŕI�(^�W8 �+N�����p��!�j�˪�U�I��}�C�����p��6����X�(*�
�x1��!�T=f� ֨3��ɽ�*<es����+���`*���Y�I��.�S�/Y:n|��(�~L�o�g�t]oA�H
E#LPA�Y��g1��0S�`O=A4C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S��!��(�V���Aj�6Q�{nvC͎B�����)�	��Ƙ����ET�:S���.8܏ ��ۆ��݋���Ƙ=���^�x�����i�]Ӕ�'�Vo�X���<FK��>I�);��K���O�dX#³�#�t�`� Dӣ�$�~�� �� ;���(Xf�F�?���܏ ��ۆ�Hlk�O3#~%w7���� *S��q�@�G�׊��.�E�� �GM;�n�a���N�sI�����F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)XC"Ɔ�;��X�
d�����d'�Z����W��M�1����?�#x8�U=�z��!�$Z��D蹯��Q� ���K�͎�U'":�L��,'�vg	?Kʩ���V]��ꘔ����	U�ݘ�=
x����}�7���kd����c�#�^���������Oz�}�F�s����G�Jct=L_ �^&��=�D蹯��Q� ���K�͎�U'":�)'Sj�~	?Kʩ���V]��ꘔ������Ci��0x����}�7���kd����c�;8*�k{T������Oz�}�F�s����G�Jct=L_ �c��M�{�D蹯��Q� ���K�͎�U'":�P�'Ϊ��	?Kʩ���V]��ꘔ����U��Fȩ�0����G�J��+��dŇN��!,YZ͆ˎ��F0k����D蹯��Q� ���K�͎�U'":�h"J���D.nxԆ&{2��Q��>֠�V�e�w�_�������G���H����$K��;��l�q���	�<���J&4L��.
��ORPB$�'�%�d���h"J���D.nxԆ&{2��Q��>֠��֋�m}]d_�������G���H����$K��;��l�q���	�<���J&4L��.
��Sc�W��%�d���h"J���D.nxԆ&{2��Q��>֠سߦ�r� i_�������G���H����$K��;��l�q���	�<���J&4L��.
��Y�iTL�둭%�d���h"J���D.nxԆ&{2��Q��>֠؇	�����_�������G���H����$K��;��l�q���	�<���J&4L��.
��q�@�+�8�%�d���h"J���D.nxԆ&{2��Q��>֠ظ�T����2_�������G���H����$K��;��l�q���	�<���J&4L��.
���9|����%�d���h"J���D.nxԆ&{2��Q��>֠�2ɂ�O�W�&x�Y�\"�ʽ;a���	�܉v��&���f���5<Im��pX(5`��q?;dh.m�14=*�D��|F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�YZ͆ˎ��~ُ��&y�.��P��D��y;W��4D<E��r;�q�C6�iM��t��[�y�i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q��H��ڟ-�ź��Z&�W�57r�<�܌��:nL�:���j`rc�d�I��ͺ����d��X��[��Ƹx���]L�E��讛 ��1�QX�k����?�ӝ����������Y ���Z&�W�B�$}�2�R���j`rc���i`��ZPL�����Y�ہ	��H���3�8�G45Z�)���=��͆����7�ž�c!J9��ӝ�����%W��G����Z&�W�B�$}�2�R���j`rc�S8Cߺ�_�PL����"TȔ��H���3�8�G45Z�)���=����t1�O���c!J9��ӝ����ܼu�"K���Z&�W�B�$}�2�R���j`rc���ˤ��PL����@�f`V�rH���3�8�G45Z�)���=����[��+t��c!J9��ӝ������P��&���Z&�W�B�$}�2�R���j`rc����$,�jPL�����v���:��H���3�8�G45Z�)���=��͵%�HW�����c!J9��ӝ�����)�A����Z&�W�B�$}�2�R���j`rc�-��hsPL������>8�2H���3�8�G45Z�)���=����|g�;Mվ�c!J9��ӝ�������7^d4�D.nxԯ�1����I��$k����xCY�R���r�m���]^�n,�Ӣ�8��Uu�B�5��$[q���L�q�����/ �y=�UU���ɖY׎�0C���>MX�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�T�N�:Y�?�v�R}ky�f˺���i�H���<��sшe>6{t�YU�f$}�xNU?�Ρe������F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)X�A)�^U�V�*�mZ4l�5cgE� �K[Γ��.L?cz�\��͢�����*j<g��"Y~:�,�2��ɖX�Mةm7���Q;�{@�EmN�
�I���*� �8z0��SҪ�X�&��%.v���+d)wq�֢��G�Q;�{@�Em�b[�l:�]0;�G�	�M��)�atBҷ��c A�[f�矑��ӆ�澮/�žC���U�8�sl�Z)^��_�����±�u<@B�Q;�{@�Em{E�6��h#A�Y��g1��0�����n�0�0��V$P��
����P댠�ܱt��oQɽ�*<e��u<@B�Q;�{@�Em�H
E#LPA�Y��gSE⫄ 2}�js���J�b�T��	ɽ�*<eúU��
���>��3uM�3pI^C�����p�����S���$e��!޷-�E������p��@9_@�R4r��O�u��N:�r�C
�V[��+�r��y����Ɔ��"C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S��)`�"���!�yC��Gc�>MFD']4�7[ğ�ka3�������kmi�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q��H��ڟ-�ź��Z&�W�57r�<�܌��!L�S����w�A�f5�*N�sv�Hn/��Be�5E�k&�r��D�l��V�,xX�u�\�Ǡ<�H��Ms��ٝ���R�W��%	A=A +'4M���/v`S^!�������D�j�)3�z���q�0��ޛfe�^C�ɽ�*<e��CǺvr���V~��0Y�P��j�H����޶(:�+�r��y�wp���	JПE�[5ɽ�*<e����
�S%iv��^����؅�LF靁�Dr�WO,!��ߋ�%�?ҦR)�oPj������~����� ���OT��:.�_ݕ�0��t!h����B���	C^�1��g�eGY��J�hu:׈S�y1bdY�D�_o��u��5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^����
�S%iv��[۪c�;���E���u�_k�=�9��+����� �}�V3����_Ai�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q�ݕ"Uy��\�V�W�v#@CH5x�`{ѕ5��l)Ȟ 胨RJПE�[5��}Gδ�-��$Q����x���]L�E��[�_�B�;�k%e\�]���tU��ɽ�*<e	?v��BR�!�	=o��R;���GN���-�8w��8t���&Nꊓ�H��䅓�g �����i88��C�3���&%�ޛfe�^C�ɽ�*<e�ӝ����vk�q嚤�L/D�%mun'(��۾/����p��Rg�9��q^�(	z��NyE,��zNh[��6����	?v��BR�|\8��>/%�������P�7ٝGy�u:׈S�yB,���m��I4������i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q�����4zm�rR��"9�I��G5)�EҀ&*����1`��sr�%�����ig���`�7L5������7�t×,3a[���ʩ�|��+��pb5�R-��	p��*�Q#B������g�XC�����M� 6%����fB4/���8\kB,����I�oPh�c��9�8Ɯ4B�PZ���]�N�� #�z�F��V(�����{N�������"-�o��
�VE�n񂰤5��:0�*�D��|F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�E��7ۅ��1��9MVqYu�ҧ�T��T�����Zm�`���j��r��O�u�H���w�b
B���^���ΦsH�Լ=�/r���m�{�e�,���WXe�]��%�0H��:����3��Υ�l����s{r@�w)�F��V(�Hy�zN�tf�1��eY`���?	�*����1`�g��+�`��X�s�J�A)�^U�#\d�^�,aΨ8��Z�D���k4�?�Vl��nE�"q��L��N�8W��O�pٺe�E��7ۅ��1��9MVq~#�m�Kqa�T��T�����Zm�`���j��r��O�u����(O
B���^���ΦsH�Լ=�/r���͓��Υ�l����s{r@�w)�F��V(��U��N�]�"8�q�R�-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�)V ٥�Dk���f�V&n����WE�"q��S�A�����9�$5<���o��K�!�@M\{�m�d��K��}�}�YZ͆ˎ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��(�'D��P������@�1�x0Yc&�r��E�"q��2�>��1���fC��F��V(��_�}d������pr��O�u�Ǫh5��P�#\d�^�,p�wV�����/�����=�/r��˿���O�^#\d�^�,�,�AA8����/�����=�/r��HU����<#\d�^�,G'+4/�\���/�����=�/r��ݺx0H
l7#\d�^�,N�Q���z���/�����=�/r����u �z�#\d�^�,P�{%������/�����=�/r��|`6S�Y�3�២x �ti�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q�݊����F2]�J8�F2]�J8�F2]�J8�F2]�J8�$�䠢O)X�A)�^U����ߓp
�	��Y��=�/r��U<�u��p�+����5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^�����qϏ�u������ZF�i��%ƨ��-�H��#��HP87ξkZ�x�'��� ���O�-�*ǻ�F�k-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��D�[m�m7���!L�]j`▘9�����V����n-�{ѕ5��l)Ȟ 胨RJПE�[5��}Gδ�-rE%R�m�O@����8T�'uw@�|��ʸhP�&Nꊓ�HU877�P�����tWɬ�l��a3#��ׂ���^*��3p~p�sQl|LF}l�.���C�3<Q��A�"Uy��\=�B��YX�>� =&d8�&��F�g���΃X��ߔG�=��C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S�ɽ�*<e��i�a/�ͷ�@�����X�eie�ȏM��8�kw�zi��sgF��G�y��_�2�Vk�'r-���E�5���(��yo�lC��m嗫�-�C�}N	2�8$���Fh��ro����n��r��<�H��Qh7�i ��i�7�;��ɽ�*<e�5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^p����N�\WjH�r�a�*�����BR�����H��z�zG�j��ґ]]���[����"�'��� d��:�cp����Nk{�nq�E�m<�z�]�}l�.����_o��u������iPt����f�\�}����u!i�l��vGU�|-W�>���D��a�DzjڢX#��<�����j`rc����.�HX�����q�E����mV����� A�[f�矑��ӆ�澮/�žC���U�8�s��c��d6VG�X�y�k[|�nRw,W�!Yn��R��_F��x��^�,�NN�F�2�pھi��͗
�m���B�R���	0Y�P���q�OO�����Ɔ��"C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S�-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�)V ٥�Dk\��kc��x�>r3�$%�5����fF2]�J8�F2]�J8�F2]�J8�F2]�J8�	C7��3�^C��ଡ଼�F2]�J8�F2]�J8�F2]�J8�F2]�J8�~�&T�S�YZ͆ˎ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��� �z F73�Z��gJb%�+�T\�28���T�k���E��C�>�_{��h���YZ͆ˎ����j����Y���Rͱ!���n�=F�
�!��)�^�ZP� mgT*�ɷ�U��8PK�XvV����r|⥫��aw����2
�t)��:>��`K^�
��VrL۪w�IbGZ)]�u��̖���u����n%D3�K��"rj�Q{��%߱��_4��X�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8�T�N�:Y�?�
���ji�:�1���-�d��\�Z�E��7ۅ���0k���ء�B�N���:nL�:���j`rc��kwu�p�w��ՌAvɽ�*<eɽ�*<eɽ�*<e�.U�[�x��Vh��;ko��ܾT#o*�L!�b��i��<�a�]�C�ﮮ���nr��<��lC��We���)e�������O��^�����	Q}.��LvԱۣq]s����'L�%'�vH�`��1�^��ש��i��@�blP�1��@\���˺�1UcjoAh�q?��y��?�$���X�Eg2�������y��ǋ2�x�Jf�q�����/ �-(�E�WȺ�����zt�](HA�6��i�S�����VM��*�a��߫;�T	�s�Gj�=�@����v�?xV���qA}��/G)�u��A��Y���t6��y��!q����`'�r�5X��,�M,�	��rɽ�*<eɽ�*<eɽ�*<eYZ͆ˎ�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8��� �z F7i�ܛ�|�F2]�J8�F2]�J8�F2]�J8�F2]�J8�����q����q26~ mgT*��o�Y�pl�'f�1!5:i���2Z����$"���h��-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�)V ٥�DkX�1�{��F2]�J8�F2]�J8�F2]�J8�F2]�J8���O��[k�����Q���Ɛ�sg��<�#Z�a�0��� �?c�5s@]?�/9
��阺����Q�	����9|�<�#Z�a�0��� �?c�5s@]?����4��t�����Q����5#����<�#Z�a�0��� �?c�5s@]?Z&ÓeȺ����Q����
��Q�<�#Z�a�0��� �?c�5s@]?J�'�B�����Q��~*&��.�<�#Z�a�0��� �?c�5s@]?��{��u������Q���(������<�#Z�a�0��� �?c�5s@]?�� ��d�����Q��)�Əƚ�<�#Z�a�0��� �?c�5s@]?�,��e������Q���z4#R
�<�#Z�a�0��� �?c�5s@]?�5�D"�4�����Q�g\;��Q���<�#Z�a�0��� �?c�5s@]?B�͝V6�����Q�]cA\=�)�<�#Z�a�0��� �?c�5s@]?W�/�S�ۺ����Q��;��,EDx����s����.�NH�*�����ɇ�ԉ���(�[�v��m$���Q
j���g���>�u=��&���?� TJ�a�i���Cf]����L��j���&��N����]Q�������r�K�+���􈂙��q�EĄ�#���K,V[d-oO�8NZ���} 7uh��F3�@rr8�?@�bZ���,��}xvI0%�����r�m���nhs;J6�@rr8�?@�bZ���,��}�c3-r\�s��r�m���1�o�5+��@rr8�?@�bZ���,��}�mR�b���r�m��͘�F"��d�@rr8�?@�bZ���,��}큵*: ;��r�m��͹Z�E�I�@rr8�?@�bZ���,��}uUbD�����r�m����y�H�6��@rr8�?@�bZ���,��}l�o���.��r�m���$�F���@rr8�?@�bZ���,��}YbՀ9 ����r�m���[��mB=�@rr8�?@�bZ���,��}����R����r�m���d��8�X�@rr8�?@�bZ���,��}����ΥmD��r�m���=|���w�@rr8�?@�bZ���,��}y����i��r�m��͏��la@:� �������!����7n�8kǪL���R��c!J9�pH[��V����{Y� N�/����2Pʍ�P֠��`�2[TS@9��-��v��,��-��KC�F2]�J8�F2]�J8�F2]�J8�F2]�J8�F2]�J8�)V ٥�Dk���� 1�$��;�P��jBC������F2]�J8�F2]�J8�F2]�J8�F2]�J8����T%�g'��^/a�m�ժ����� ���rܬ`T��8����c���`iF�-��yN�F�8I7uh��F3�����d<�������|Gb��f	>����̓4����?5V �y�l��,t	 kp(���&b���z&�Y����X�y4{j�}pH[��V�	/wx�ۻ���F����OG����`�K�am@���JyĥQGi
��Cj��[�j����6VN�9�g�'m�L������'�z�XQ�,������oN��m�B���z%s��:˃�6��RbD:�I�M�}��Pj���"�q����9��p���7/'��������ߢ���&��!Q]��ھ�>j}�!�(I�J��'�U��!��/Ϫg���4`՝�^/a�hТ�z�I}� ���rܬ`T��{/U Qz�<���ae`�yN�F�8I�Z�E�I�����d<�������2Nf*v�"�����̓4����?5V �y�l�� W���Ib(���&b��,mɺ�ǴY����X��2��pH[��V���(�4�1���F���1�׷))Y��K�am@���JyĥQGi
��Cj�l�Q(����6VN�9� �:+|<�����T��N�,�,�����.��b��Lm�B���gϥ�\�� ˃�6��RbD:�I�M�}��Pjw����/���9��ͮ�s���6'���x�9:��i��&��!Q]8p�!���!�(I�J��'�U����3\�����4`՝�^/a�j����4=�� ���rܬ`T������#z;�1��yN�F�8Id��8�X�����d<�������1J9S�~������̓4����?5V �y�l��Hм&�Su(���&bF �<�*�Y����X��\��pH[��V���D8QXzȓ�F����seFxG&��K�am@���JyĥQGi
��Cj�LaQ�y��9�t& ҿà��s�'���ff�:?�~ȅ�J�_��!)k0�[�����d<������Ԡ���@a�V8��+ Z&�s�����u��_a�#-�s�S��6VN�9�`Mg������D���ob ��5R�I��&��!Q]�x���KG5�td'�44�Ik�PCZ�\:�(����̓4k�N*�%��Û�ff�����g�@P�c��9�OఓG~��砽���d<�
a�E��z����v��{�^�W�n�����&-�G�l����`1��������{9�\4�"�ѫyt,A�~ړ��4E�{�^�'V�W,9�{M���S�w�s@�����4�
��������iq�f��>��D����N�,9�{M���)_d<�cYb�'����4�È}����Hc�;�Y^�U=���8��u��w��湬��>n.r�P�S��И]h����,��D�se��L���Ӡ��B:l��9q؟��?��6���꨽�I0B�O�F��֕pR�Lʉ/[¶���`���c��� �	[�w:���ע��������t��$:ԑ"�C�#1���a��0�[��z����jcbb_�B�,��y8f���B6Km���'�5uEq_�<|7.�n�B�D���|�w��M{�˦��w1_#Ǚ��R�����'c.�	?0-� ����Jv�T�`���LZu��,��m#u01gHg)%�RPz
2����
�7`�	�6��o�y!��;��od<~��Og6i���H����I��	n�2�Y�RoѼ5T�g�'y{�I��y3AL�����~ָ���}R�|��`iX��-m$�V��o����W�d��\A�\��B�1U�<`<�a[��6����J�
��\�O����7�X5/�)1@U����݋�Ǹ�
���������h�>K	�K�7	�j����m%p7m�R���|"ÝW�qe�
��Wi�5��������̹�"�j��;�kԐH`�Q�;sXf�D�V�²z<rt�����}3�Wџ5)l`�AG�0����{d�����V�²z<rt�����-Q�*����'��.�X�O��]vMEZ1�*�=m?!~�H�^U_�>�5?�;�|���0�*G �l8��xȺ���jd��3��W�<�)>�YG �l8�永�`�R꾯a�F�zM�����3��6�4�#�ՙ6Nk%-�ư�=���g���f+�ph9!�4�hԚԾ3��R
y�h�ᕑxpu��8B`}������ɽ�*<eɽ�*<eɽ�*<e�VJUT���!�vh!T	�B迸Ψ�ɽ�*<eɽ�*<eɽ�*<e�cǭ����(��^o�ɽ�*<eɽ�*<eɽ�*<e:j���+�Xq��hH�ɽ�*<eɽ�*<eɽ�*<e�&�|�D��_���V��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�&Z6[�f�UgYavɽ�*<eɽ�*<eɽ�*<eZC���O��~bj�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eA�w��usR�fs!_ɽ�*<eɽ�*<eɽ�*<e`�!ܒ������N���6�8��'�^���:4���7�m��p~A9����W�Z��J�j��1H�f{��~��Wɽ�*<e	�������~��Wإ�'C8�/xQP�?@����㭊x�.�^<�
:�vS+ё@OXSf��D�5�j���ɽ�*<e?���Y����_���2"\�>����$�"`��x��$�?5��vʁ��H�?i�����Z�`õ�|�M�ʟ��k �S��t�6�Z��Ѣ��Y�8�����Q�t���@��!���,TV�J�U�d]7jȫ������Y�](�����������Q��s�8RSJ�&&��k��Y}���ǈ��� *B�Ե�5���bl��"Uy��\�V�W�v#@CH5x�`|�L��y�w�&Z6[��խ|��e�k���,(n���M���Nl1p�N&�]����i{ޝ��i��':y����g���wp���	�?�rm���(����i{ޝ��i��':y�{����e�m5�1g$��{��t6��_0(������9n;NǕl1CQ���!��4�,@hp��Ԁ�F�Y���~N�� ���}���bU���z~@�U��t����{����f�2_B@�~%.DI���:��t�%2����TW�lZC���,<�r���+9}�t����{����f�2_B@:P��dS	nT��e�&��F]�J�������	U�֝�%��L�f��iq]��
�k���_=������Y�"�WZ9���u\�a݀P�!s�,�	���Π�އ�Fs��s+s�ߥ�x��!6���f����!Lؒ&�bL�.��. ����lB��,zyj���0_��A�\��B�o�����'�)��<L}ڈ�����dn'y&���3��ͨL���K��a9q;���]��e�G<���ߤ#� ����2W�rB�������i0��|"ÝW}�utiO����+�%�Q)=d���E@�׺�F�b3��5�э1��!S�)����qӬ�\ԗ�fd�5�\� �zņ�m]1��F�^v�'-�cb�S���mheˣ����ܯN�ՃuL�7d̈w�U���YEL8��L�Y���ay\�n ���J?|��'����A�as��MF�R�i ��֔��a�uP�M�z�ڽS7��v�����
����%�z�M	!���=��ϝ�p:�\���YV��������m\R��Ey�>�t�Jд��߿Kv���������0���L��J���n�+cb�p�W�f�ܑk���g+��jj�h��#B�`b��-����6�cW�n2L�CA�A~R��72���؛��}s0�0�Q�����6�cW�n2dꜱ+�	��������"!f5@fF� >����� Y����p��x����f��e�*�=o�ZL9���D�>'TP%0MA��x�<:?w��J8�q9���D�>'TP%0MA�Q�S��-Ye@�M�����a��	P���Z����5���\+��b�ε�,Y�^e[��z��I-��c���A��G��x�]�ͻlU��]@x0�z�ɽ�*<eɽ�*<eɽ�*<e�VJUT���!�vh!T	�B迸Ψ�ɽ�*<eɽ�*<eɽ�*<e���7	��lb�`i�Iɽ�*<eɽ�*<eɽ�*<eܞ�P�c]��c�u�h[�����p��ɽ�*<eɽ�*<eɽ�*<e>"��;a��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�.��W�����p��ɽ�*<eɽ�*<eɽ�*<e��`V�;�.�]� ��)!ɽ�*<eɽ�*<eɽ�*<e0������ޟ:k���ɽ�*<eɽ�*<eɽ�*<eɽ�*<eY��>t���!x"�#��ɽ�*<eɽ�*<eɽ�*<e]�P�.�F_���V��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e/���?������p��ɽ�*<eɽ�*<e~M3Y����)�y��g�i�py�h�*`�8�Pϟn�Cb���A|�eP�[N�b��AB�O�aS�O�. ���\�I;�����l3!���p��S	��ػN0B��wo�	h�[ܞ�P�c]��:sv�]�9�ψ���ɽ�*<eV���X�f�9�ψ���ɽ�*<e7��� h�4b�]��C5����_k`ɽ�*<e���@=n�9�ψ���Hpm��A�,h9IO��^b�����E]�d���B�ɽ�*<e��]��.58����Kċ����$5�g���D�E�? ^����vʁ��H9q�[[��	��l����ZV�����/��Bg����U�酎�P�#�L����+��ȉ�/���?��z5ߘ�严%�;�"�,��
�L���-,�Deϑ���O�ۚ�(�,<h�$�5:���p���D.����LJ�ڤ���$ys2��4�>I��\����Br��pE��7�αNa����G���R�ʹXr�I,N��o+m��Fo�ly+�7��	t�nQ���
����+(M�e~�MI�䕟�ɽ�*<e��YqF��^����.?��&Nꊓ�Ho�
�0�C��_�av"#x^�4�4s��7�+��s�a2궼<<mP��7�ھi��͗
�^��"�6�t�V�,�i���!�)�ny�Qu�3���_0(������лV�|�®�O���}U�b,� �%��Bg����)�D��c}��Pj�/��5ı��>�j*�r����A��mt�[���{9�����b}V�yt,A�~ړ��4E�{�^�'V�W,9�{M���S�w�s@�����4�
��������iq�f��>��D����N�,9�{M���)_d<�cYb�'����4�È}����Hc�;�Y^�U=���8��u��w��湬��>n.r�P�S��И]h����,��D�se��L���Ӡ��B:l��9q؟��?��6���꨽�I0B�O�F��֕pR�Lʉ/[¶���`���c��� �	[�w:���ע��������t��$:ԑ"�C�#1���a��0�[��z����jcbb_�B�,��y8f���B6Km���'�5uEq_�<|7.�n�B�D���|�w��M{�˦��w1_#Ǚ��R�����'c.�	?0-� ����Jv�T�`���LZu��,��m#u01gHg)%�RPz
2����
�7`�	�6��o�y!��;��od<~��Og6i���H����I��	n�2�Y�RoѼ5T�g�'y{�I��y3AL�����~ָ���}R�|��`iX��-m$�V��o����W�d��\A�\��B�1U�<`<�a[��6����J�
��\�O����7�X5/�)1@U����݋�Ǹ�
���������h�>K	�K�7	�j����m%p7m�R���|"ÝW�qe�
��Wi�5��������̹�"�j��;�kԐH`�Q�;sXf�D�V�²z<rt�����}3�Wџ5)l`�AG�0����{d�����V�²z<rt�����-Q�*����'��.�X�O��]vMEZ1�*�=m?!~�H�^U_�>�5?�;�|���0�*G �l8��xȺ���jd��3��W�<�)>�YG �l8�永�`�R꾯a�F�zM�����3��6�4�#�ՙ6Nk%-�ư�=���g���f+�ph9!�4�hԚԾ3��R
y�h��~��=����8B`}������ɽ�*<eɽ�*<eɽ�*<e�VJUT���!�vh!T	�B迸Ψ�ɽ�*<eɽ�*<eɽ�*<e�cǭ����(��^o�ɽ�*<eɽ�*<eɽ�*<e:j���+�Xq��hH�ɽ�*<eɽ�*<eɽ�*<e�&�|�D��_���V��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�&Z6[�f�UgYavɽ�*<eɽ�*<eɽ�*<eZC���O��~bj�ɽ�*<eɽ�*<eɽ�*<eɽ�*<eA�w��usR�fs!_ɽ�*<eɽ�*<eɽ�*<e`�!ܒ������N���6�8��'�^���:4���7�m��p~A9����W�Z��J�j��1H�f{��~��Wɽ�*<e	�������~��W�@P�/xQP�?@����㭊x�.�^<�
:�vS+ё@OXSf��D�5�j���ɽ�*<e?���Y����_���2��i5=9����$�"`��x��$�?5��vʁ��H�@�c���Z�`õ�|�M�ʟ��k �S��t�6�Z��Ѣ��Y�8�����Q�t���@��!���,TV�J�U�d]7jȫ������Y�](�����������Q��s�8RSJ�&&��k�P&n�(��L�ǈ��� *B�Ե�5���bl��"Uy��\�V�W�v#@CH5x�`|�L��y�w�&Z6[��խ|��e�k���,(n���M���Nl1p�N&�]����i{ޝ��i��':y����g���wp���	�?�rm���(����i{ޝ��i��':y�{����e�m5�1g$��{��t6��_0(������9n;NǕl1CQ���!��4�,@hp��Ԁ�F�Y���~N�VB������}���bU���z~@�U��t����{����f�2_B@�~%.DI���:��t�%2����TW�lZC���,<�r���+9}�t����{����f�2_B@:P��dS	nT��e�&��F]�J�������	U�֝�%��L�f��iq]��
�k���_=������Y�"�WZ9���u\�a݀P�!s�,�	���Π�އ�Fs��s+s�ߥ�x��!6���f����!Lؒ&�bL�.��. ����lB��,zyj���0_��A�\��B�o�����'�)��<L}ڈ�����dn'y&���3��ͨL���K��a9q;���]��e�G<���ߤ#� ����2W�rB�������i0��|"ÝW}�utiO����+�%�Q)=d���E@�׺�F�b3��5�э1��!S�)����qӬ�\ԗ�fd�5�\� �zņ�m]1��F�^v�'-�cb�S���mheˣ����ܯN�ՃuL�7d̈w�U���YEL8��L�Y���ay\�n ���J?|��'����A�as��MF�R�i ��֔��a�uP�M�z�ڽS7��v�����
����%�z�M	!���=��ϝ�p:�\���YV��������m\R��Ey�>�t�Jд��߿Kv���������0���L��J���n�+cb�p�W�f�ܑk���g+��jj�h��#B�`b��-����6�cW�n2L�CA�A~R��72���؛��}s0�0�Q�����6�cW�n2dꜱ+�	��������"!f5@fF� >����� Y����p��x����f��e�*�=o�ZL9���D�>'TP%0MA��x�<:?w��J8�q9���D�>'TP%0MA�Q�S��-Ye@�M�����a��	P���Z����5���\+��b�ε�,Y�^e[��z��I-��c���A��t^��λq f�&��p��ɽ�*<eɽ�*<eɽ�*<eɽ�*<e(���٤r�!x"�#��ɽ�*<eɽ�*<eɽ�*<eL�r��NBs郝���ɽ�*<eɽ�*<eɽ�*<eɽ�*<e���.���ɽ�*<eɽ�*<eɽ�*<eɽ�*<e�� �X������p��ɽ�*<eɽ�*<eɽ�*<e`ύ���#��I�~�	ɽ�*<eɽ�*<eɽ�*<e,4���?w�<y���$�B迸Ψ�ɽ�*<eɽ�*<eɽ�*<e��ky�-��'(f9��ɽ�*<eɽ�*<eɽ�*<eL��]�1�A|�eP�[N�b��AB�O�aS�O�. ���\�I;�����l3!���p��S	��ػN0B��wo�	h�[���r�<ػN0B��+b�6����O��xx����W��\�I;���ɽ�*<e�&Z6[��u�ᐣ�ɽ�*<e���r�<������]���>�c��T�F�v�N����P��#�L��׸
������s�8RSJ7�\ �9~d;#R��ot���X�N�`?=>YJ�l�EX�F���$�_K�Y�nX�M��h�o�T��0��(/�� ��U�L>YJ�l�E���T��Ќv���t����%��8�2��4�>I��\����BfbeB܃'JFP������.
�_F��D��k��-�]d���)%��b0�4�v	;o�`V�f�BO�
�����p��V�e�><��P%ɽ�*<e3\�!ќ��M�=�8��ŕI�(^�F��Ư@��
&�ɽ�*<e3\�!ќ���5i��̕��0����Z�`õ�%o�g�~V�[еP�����Q�=w�,lD��d6��`��y��M�&������Uj����}�����&j:o�$�T���]��q`=��ϝ�p:��
D��H���/T� ���\����q�:�Ʈ�<#JZ,�:�Ek=��ϝ�p:��
D��H7����{�ƥUuh��V�g5D�l��9q�X�:׮�{k��kx6�j��"�yL�x���Ys�}�q��?Xٵ��5�,����F]�J�������	UQQ*rb���f̟�zǎQe�[D���bc+Ji �8s����6e���%���2"��
��4N;L�Oc]���2��sbK���P@Q|b�`�/^�:���;⑤���a,�"�빱x�Q<�^eg��ɂ����c_�o� x/���z�����i���KDh�D;&��'���b���Ly�|y�ި���6�ʈ����I;��?d�o h�o�c�N���Īö�{T��qɮ��B���(���%��|`ଽ��p�N_�qe�
��bS�����"�N�?�����LV���:Wp<!���I��d�>�r=D�9�)�Ί#|�Ӏm��!Q	s>R=��@A��\��G	�#1
 H��D�����e�mu���H��H�
:��p��؋9i��������a:�#�f"��]b9�`�u�ת���A �Ы���VI#�1z���x�q��Ǝ�b\[��½�#��$̆���5��0�F�P$��Vڸ4��| ���Xj��)�*��e/6�5��0�򐹸���9��/BƷ?�yN��d3M6�YLQg8l&�cψ5���Jt��ٍ��WF��洴�/BƷ?�yN��d3M6�˨
�c�pp&�\Գ�cl&��l@��1�9�vd&DzR�5'(�H,[As�M�Z���FB�qxj3T�zm�Jw��8ht]ٽ�x���FB�qxj3T�zZ����(�
-İx��s�JV�^��_@�Y�x��g)^�՘&7(� J)�͕[����oz)���ʠ��6�x�A-��b=��K�X���hs������p��ɽ�*<eɽ�*<eɽ�*<e) uN)BQ��7�����ɽ�*<eɽ�*<eɽ�*<e���7	��lb�`i�Iɽ�*<eɽ�*<eɽ�*<e�%��IC�KS�E`�jdɽ�*<eɽ�*<eɽ�*<eɽ�*<eT#@�GNɽ�*<eɽ�*<eɽ�*<e��_��l���]V&a;Bɽ�*<eɽ�*<eɽ�*<e�����>xs1�|�ɽ�*<eɽ�*<eɽ�*<e"7�!ne*5^|��]`�f�UgYavɽ�*<eɽ�*<eɽ�*<e�s��"�w�[g�Ʊ�]ɽ�*<eɽ�*<eɽ�*<e���&B��29'�ɽ�*<eɽ�*<eɽ�*<eɽ�*<e/���?������p��ɽ�*<eɽ�*<e"4�R��׾υ��.�ɜ�S��җ�f$�v�*[��	��l���W<:K�k����Gv_^���_�F�?�C9�Ru�:\_�k�:a���i ��
��R'9�ψ���ɽ�*<e�%��IC�KQ���h��~��Wɽ�*<e	�������~��Wɽ�*<e`ύ���#M���nz�~.�^<�
:�"7�!ne*5[�q5�s���~��W�k����Gv�M��GW%}���!����Zɽ�*<e�c��_��P���������.rݸ�mnp i�ij����ȵ��t����I�e�g���A�#�L��׸
������s�8RSJ|�Jv@�f��_��Tㄽot���X�N�`?=>YJ�l�EX�F���$�_K�Y�nX�M��h�o�T��0��(/�� ��U�L>YJ�l�E���T��Ќv���t����%��8�2��4�>I��\����Br��pE��7�αNa����G���R�ʹXr�I,N��o+m��Fo�ly+�7��	t�nQ���
����+(M�e~�MI�䕟�ɽ�*<e��YqF��^����.?��&Nꊓ�Ho�
�0�C��_�av"#x^�4�4s��7�+��s�a2궼<<mP��7�ھi��͗
�^��"�6�t�V�,�i���!�)۞�:"�d��{Vent�Ŏǣ�[Ƹ5��X�p zpM���:".�~�bW\-k�*���fv>YJ�l�E7�.봹�r��>���_ I]f�Yj}Rk!��ʛ�uK!b�b*A��